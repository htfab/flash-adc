magic
tech sky130A
magscale 1 2
timestamp 1713341356
<< metal2 >>
rect 8556 37992 8616 38001
rect 8556 37923 8616 37932
rect 8924 37992 8984 38001
rect 8924 37923 8984 37932
rect 9292 37992 9352 38001
rect 9292 37923 9352 37932
rect 9660 37992 9720 38001
rect 9660 37923 9720 37932
rect 10028 37992 10088 38001
rect 10028 37923 10088 37932
rect 10396 37992 10456 38001
rect 10396 37923 10456 37932
rect 10764 37992 10824 38001
rect 10764 37923 10824 37932
rect 11132 37992 11192 38001
rect 11132 37923 11192 37932
rect 11500 37992 11560 38001
rect 11500 37923 11560 37932
rect 11868 37992 11928 38001
rect 11868 37923 11928 37932
rect 12236 37992 12296 38001
rect 12236 37923 12296 37932
rect 12604 37992 12664 38001
rect 12604 37923 12664 37932
rect 12972 37992 13032 38001
rect 12972 37923 13032 37932
rect 13340 37992 13400 38001
rect 13340 37923 13400 37932
rect 13708 37992 13768 38001
rect 13708 37923 13768 37932
rect 14076 37992 14136 38001
rect 14076 37923 14136 37932
rect 14444 37992 14504 38001
rect 14444 37923 14504 37932
rect 14812 37992 14872 38001
rect 14812 37923 14872 37932
rect 15180 37992 15240 38001
rect 15180 37923 15240 37932
rect 15548 37992 15608 38001
rect 15548 37923 15608 37932
rect 15916 37992 15976 38001
rect 15916 37923 15976 37932
rect 16284 37992 16344 38001
rect 16284 37923 16344 37932
rect 16652 37992 16712 38001
rect 16652 37923 16712 37932
rect 17020 37992 17080 38001
rect 17020 37923 17080 37932
rect 17388 37992 17448 38001
rect 17388 37923 17448 37932
rect 17756 37992 17816 38001
rect 17756 37923 17816 37932
rect 18124 37992 18184 38001
rect 18124 37923 18184 37932
rect 18492 37992 18552 38001
rect 18492 37923 18552 37932
rect 18860 37992 18920 38001
rect 18860 37923 18920 37932
rect 19228 37992 19288 38001
rect 19228 37923 19288 37932
rect 19596 37992 19656 38001
rect 19596 37923 19656 37932
rect 19964 37992 20024 38001
rect 19964 37923 20024 37932
rect 20332 37992 20392 38001
rect 20332 37923 20392 37932
rect 20700 37992 20760 38001
rect 20700 37923 20760 37932
rect 21068 37992 21128 38001
rect 21068 37923 21128 37932
rect 21436 37992 21496 38001
rect 21436 37923 21496 37932
rect 21804 37992 21864 38001
rect 21804 37923 21864 37932
rect 22172 37992 22232 38001
rect 22172 37923 22232 37932
rect 22540 37992 22600 38001
rect 22540 37923 22600 37932
rect 22908 37992 22968 38001
rect 22908 37923 22968 37932
rect 8558 37860 8614 37923
rect 8926 37860 8982 37923
rect 9294 37860 9350 37923
rect 9662 37860 9718 37923
rect 10030 37860 10086 37923
rect 10398 37860 10454 37923
rect 10766 37860 10822 37923
rect 11134 37860 11190 37923
rect 11502 37860 11558 37923
rect 11870 37860 11926 37923
rect 12238 37860 12294 37923
rect 12606 37860 12662 37923
rect 12974 37860 13030 37923
rect 13342 37860 13398 37923
rect 13710 37860 13766 37923
rect 14078 37860 14134 37923
rect 14446 37860 14502 37923
rect 14814 37860 14870 37923
rect 15182 37860 15238 37923
rect 15550 37860 15606 37923
rect 15918 37860 15974 37923
rect 16286 37860 16342 37923
rect 16654 37860 16710 37923
rect 17022 37860 17078 37923
rect 17390 37860 17446 37923
rect 17758 37860 17814 37923
rect 18126 37860 18182 37923
rect 18494 37860 18550 37923
rect 18862 37860 18918 37923
rect 19230 37860 19286 37923
rect 19598 37860 19654 37923
rect 19966 37860 20022 37923
rect 20334 37860 20390 37923
rect 20702 37860 20758 37923
rect 21070 37860 21126 37923
rect 21438 37860 21494 37923
rect 21806 37860 21862 37923
rect 22174 37860 22230 37923
rect 22542 37860 22598 37923
rect 22910 37860 22966 37923
rect 8650 27308 8706 31190
rect 7362 27252 8706 27308
rect 7362 26052 7419 27252
rect 9662 27108 9718 31190
rect 7682 27052 9718 27108
rect 7682 26052 7738 27052
rect 10674 26908 10730 31190
rect 11686 27308 11742 31190
rect 12698 27308 12754 31190
rect 11686 27252 11838 27308
rect 8002 26852 10730 26908
rect 8002 26053 8059 26852
rect 8002 26052 8058 26053
rect 11781 26052 11838 27252
rect 12092 27252 12754 27308
rect 12092 26052 12150 27252
rect 13710 27108 13766 31190
rect 12422 27085 13766 27108
rect 12420 27052 13766 27085
rect 12420 26052 12478 27052
rect 14722 26908 14778 31190
rect 15734 27308 15790 30948
rect 16746 27308 16802 31190
rect 15734 27252 16368 27308
rect 12732 26852 14778 26908
rect 12732 26053 12789 26852
rect 12732 26052 12788 26053
rect 16312 26052 16368 27252
rect 16632 27252 16802 27308
rect 16632 26052 16688 27252
rect 17758 27108 17814 31190
rect 16952 27052 17814 27108
rect 16952 26052 17008 27052
rect 18770 26908 18826 31190
rect 17272 26852 18826 26908
rect 19782 26908 19838 31190
rect 20794 27108 20850 31190
rect 21806 27108 21862 31190
rect 20794 27052 21218 27108
rect 19782 26852 20898 26908
rect 17272 26052 17328 26852
rect 20842 26052 20898 26852
rect 21162 26052 21218 27052
rect 21482 27052 21862 27108
rect 21482 26052 21538 27052
rect 22818 26908 22874 31190
rect 21802 26852 22874 26908
rect 21802 26052 21858 26852
rect 7369 26051 7419 26052
rect 11781 26051 11831 26052
rect 12420 26051 12470 26052
rect 16312 26051 16362 26052
rect 16953 26051 17003 26052
rect 20844 26051 20894 26052
rect 21484 26051 21534 26052
<< via2 >>
rect 8556 37932 8616 37992
rect 8924 37932 8984 37992
rect 9292 37932 9352 37992
rect 9660 37932 9720 37992
rect 10028 37932 10088 37992
rect 10396 37932 10456 37992
rect 10764 37932 10824 37992
rect 11132 37932 11192 37992
rect 11500 37932 11560 37992
rect 11868 37932 11928 37992
rect 12236 37932 12296 37992
rect 12604 37932 12664 37992
rect 12972 37932 13032 37992
rect 13340 37932 13400 37992
rect 13708 37932 13768 37992
rect 14076 37932 14136 37992
rect 14444 37932 14504 37992
rect 14812 37932 14872 37992
rect 15180 37932 15240 37992
rect 15548 37932 15608 37992
rect 15916 37932 15976 37992
rect 16284 37932 16344 37992
rect 16652 37932 16712 37992
rect 17020 37932 17080 37992
rect 17388 37932 17448 37992
rect 17756 37932 17816 37992
rect 18124 37932 18184 37992
rect 18492 37932 18552 37992
rect 18860 37932 18920 37992
rect 19228 37932 19288 37992
rect 19596 37932 19656 37992
rect 19964 37932 20024 37992
rect 20332 37932 20392 37992
rect 20700 37932 20760 37992
rect 21068 37932 21128 37992
rect 21436 37932 21496 37992
rect 21804 37932 21864 37992
rect 22172 37932 22232 37992
rect 22540 37932 22600 37992
rect 22908 37932 22968 37992
<< metal3 >>
rect 778 45142 878 45152
rect 778 44962 788 45142
rect 868 44962 878 45142
rect 778 44952 878 44962
rect 1514 45142 1614 45152
rect 1514 44962 1524 45142
rect 1604 44962 1614 45142
rect 1514 44952 1614 44962
rect 2250 45142 2350 45152
rect 2250 44962 2260 45142
rect 2340 44962 2350 45142
rect 2250 44952 2350 44962
rect 2986 45142 3086 45152
rect 2986 44962 2996 45142
rect 3076 44962 3086 45142
rect 2986 44952 3086 44962
rect 3722 45142 3822 45152
rect 3722 44962 3732 45142
rect 3812 44962 3822 45142
rect 3722 44952 3822 44962
rect 4458 45142 4558 45152
rect 4458 44962 4468 45142
rect 4548 44962 4558 45142
rect 4458 44952 4558 44962
rect 5194 45142 5294 45152
rect 5194 44962 5204 45142
rect 5284 44962 5294 45142
rect 5194 44952 5294 44962
rect 5930 45142 6030 45152
rect 5930 44962 5940 45142
rect 6020 44962 6030 45142
rect 5930 44952 6030 44962
rect 6666 45142 6766 45152
rect 6666 44962 6676 45142
rect 6756 44962 6766 45142
rect 6666 44952 6766 44962
rect 7402 45142 7502 45152
rect 7402 44962 7412 45142
rect 7492 44962 7502 45142
rect 7402 44952 7502 44962
rect 8138 45142 8238 45152
rect 8138 44962 8148 45142
rect 8228 44962 8238 45142
rect 8138 44952 8238 44962
rect 8874 45142 8974 45152
rect 8874 44962 8884 45142
rect 8964 44962 8974 45142
rect 8874 44952 8974 44962
rect 9610 45142 9710 45152
rect 9610 44962 9620 45142
rect 9700 44962 9710 45142
rect 9610 44952 9710 44962
rect 10346 45142 10446 45152
rect 10346 44962 10356 45142
rect 10436 44962 10446 45142
rect 10346 44952 10446 44962
rect 11082 45142 11182 45152
rect 11082 44962 11092 45142
rect 11172 44962 11182 45142
rect 11082 44952 11182 44962
rect 11818 45142 11918 45152
rect 11818 44962 11828 45142
rect 11908 44962 11918 45142
rect 11818 44952 11918 44962
rect 12554 45142 12654 45152
rect 12554 44962 12564 45142
rect 12644 44962 12654 45142
rect 12554 44952 12654 44962
rect 13290 45142 13390 45152
rect 13290 44962 13300 45142
rect 13380 44962 13390 45142
rect 13290 44952 13390 44962
rect 14026 45142 14126 45152
rect 14026 44962 14036 45142
rect 14116 44962 14126 45142
rect 14026 44952 14126 44962
rect 14762 45142 14862 45152
rect 14762 44962 14772 45142
rect 14852 44962 14862 45142
rect 14762 44952 14862 44962
rect 15498 45142 15598 45152
rect 15498 44962 15508 45142
rect 15588 44962 15598 45142
rect 15498 44952 15598 44962
rect 16234 45142 16334 45152
rect 16234 44962 16244 45142
rect 16324 44962 16334 45142
rect 16234 44952 16334 44962
rect 16970 45142 17070 45152
rect 16970 44962 16980 45142
rect 17060 44962 17070 45142
rect 16970 44952 17070 44962
rect 17706 45142 17806 45152
rect 17706 44962 17716 45142
rect 17796 44962 17806 45142
rect 17706 44952 17806 44962
rect 18442 45142 18542 45152
rect 18442 44962 18452 45142
rect 18532 44962 18542 45142
rect 18442 44952 18542 44962
rect 19178 45142 19278 45152
rect 19178 44962 19188 45142
rect 19268 44962 19278 45142
rect 19178 44952 19278 44962
rect 19914 45142 20014 45152
rect 19914 44962 19924 45142
rect 20004 44962 20014 45142
rect 19914 44952 20014 44962
rect 20650 45142 20750 45152
rect 20650 44962 20660 45142
rect 20740 44962 20750 45142
rect 20650 44952 20750 44962
rect 21386 45142 21486 45152
rect 21386 44962 21396 45142
rect 21476 44962 21486 45142
rect 21386 44952 21486 44962
rect 22122 45142 22222 45152
rect 22122 44962 22132 45142
rect 22212 44962 22222 45142
rect 22122 44952 22222 44962
rect 22858 45142 22958 45152
rect 22858 44962 22868 45142
rect 22948 44962 22958 45142
rect 22858 44952 22958 44962
rect 23594 45142 23694 45152
rect 23594 44962 23604 45142
rect 23684 44962 23694 45142
rect 23594 44952 23694 44962
rect 24330 45142 24430 45152
rect 24330 44962 24340 45142
rect 24420 44962 24430 45142
rect 24330 44952 24430 44962
rect 25066 45142 25166 45152
rect 25066 44962 25076 45142
rect 25156 44962 25166 45142
rect 25066 44952 25166 44962
rect 25802 45142 25902 45152
rect 25802 44962 25812 45142
rect 25892 44962 25902 45142
rect 25802 44952 25902 44962
rect 26538 45142 26638 45152
rect 26538 44962 26548 45142
rect 26628 44962 26638 45142
rect 26538 44952 26638 44962
rect 27274 45142 27374 45152
rect 27274 44962 27284 45142
rect 27364 44962 27374 45142
rect 27274 44952 27374 44962
rect 28010 45142 28110 45152
rect 28010 44962 28020 45142
rect 28100 44962 28110 45142
rect 28010 44952 28110 44962
rect 28746 45142 28846 45152
rect 28746 44962 28756 45142
rect 28836 44962 28846 45142
rect 28746 44952 28846 44962
rect 29482 45142 29582 45152
rect 29482 44962 29492 45142
rect 29572 44962 29582 45142
rect 29482 44952 29582 44962
rect 798 38190 858 44952
rect 1534 38390 1594 44952
rect 2270 38590 2330 44952
rect 3006 38790 3066 44952
rect 3742 38990 3802 44952
rect 4478 39190 4538 44952
rect 5214 39390 5274 44952
rect 5950 39590 6010 44952
rect 6686 39790 6746 44952
rect 7422 39990 7482 44952
rect 8158 40190 8218 44952
rect 8894 40390 8954 44952
rect 9630 40590 9690 44952
rect 10366 40790 10426 44952
rect 11102 40990 11162 44952
rect 11838 41190 11898 44952
rect 12574 41390 12634 44952
rect 13310 41590 13370 44952
rect 14046 41790 14106 44952
rect 14782 41990 14842 44952
rect 15518 42190 15578 44952
rect 15518 42130 15976 42190
rect 14782 41930 15608 41990
rect 14046 41730 15240 41790
rect 13310 41530 14872 41590
rect 12574 41330 14504 41390
rect 11838 41130 14136 41190
rect 11102 40930 13768 40990
rect 10366 40730 13400 40790
rect 9630 40530 13032 40590
rect 8894 40330 12664 40390
rect 8158 40130 12296 40190
rect 7422 39930 11928 39990
rect 6686 39730 11560 39790
rect 5950 39530 11192 39590
rect 5214 39330 10824 39390
rect 4478 39130 10456 39190
rect 3742 38930 10088 38990
rect 3006 38730 9720 38790
rect 2270 38530 9352 38590
rect 1534 38330 8984 38390
rect 798 38130 8616 38190
rect 8556 38038 8616 38130
rect 8924 38038 8984 38330
rect 9292 38038 9352 38530
rect 9660 38038 9720 38730
rect 10028 38038 10088 38930
rect 10396 38038 10456 39130
rect 10764 38038 10824 39330
rect 11132 38038 11192 39530
rect 11500 38038 11560 39730
rect 11868 38038 11928 39930
rect 12236 38038 12296 40130
rect 12604 38038 12664 40330
rect 12972 38038 13032 40530
rect 13340 38038 13400 40730
rect 13708 38038 13768 40930
rect 14076 38038 14136 41130
rect 14444 38038 14504 41330
rect 14812 38038 14872 41530
rect 15180 38038 15240 41730
rect 15548 38038 15608 41930
rect 15916 38038 15976 42130
rect 16254 38190 16314 44952
rect 16990 41590 17050 44952
rect 16652 41530 17050 41590
rect 16254 38130 16344 38190
rect 16284 38038 16344 38130
rect 16652 38038 16712 41530
rect 17726 41390 17786 44952
rect 17020 41330 17786 41390
rect 17020 38038 17080 41330
rect 18462 41190 18522 44952
rect 17388 41130 18522 41190
rect 17388 38038 17448 41130
rect 19198 40990 19258 44952
rect 17756 40930 19258 40990
rect 17756 38038 17816 40930
rect 19934 40790 19994 44952
rect 18124 40730 19994 40790
rect 18124 38038 18184 40730
rect 20670 40590 20730 44952
rect 18492 40530 20730 40590
rect 18492 38038 18552 40530
rect 21406 40390 21466 44952
rect 18860 40330 21466 40390
rect 18860 38038 18920 40330
rect 22142 40190 22202 44952
rect 19228 40130 22202 40190
rect 19228 38038 19288 40130
rect 22878 39990 22938 44952
rect 19596 39930 22938 39990
rect 19596 38038 19656 39930
rect 23614 39790 23674 44952
rect 19964 39730 23674 39790
rect 19964 38038 20024 39730
rect 24350 39590 24410 44952
rect 20332 39530 24410 39590
rect 20332 38038 20392 39530
rect 25086 39390 25146 44952
rect 20700 39330 25146 39390
rect 20700 38038 20760 39330
rect 25822 39190 25882 44952
rect 21068 39130 25882 39190
rect 21068 38038 21128 39130
rect 26558 38990 26618 44952
rect 21436 38930 26618 38990
rect 21436 38038 21496 38930
rect 27294 38790 27354 44952
rect 21804 38730 27354 38790
rect 21804 38038 21864 38730
rect 28030 38590 28090 44952
rect 22170 38530 28090 38590
rect 22172 38038 22232 38530
rect 28766 38390 28826 44952
rect 22540 38330 28826 38390
rect 22540 38038 22600 38330
rect 29502 38190 29562 44952
rect 22908 38130 29562 38190
rect 22908 38038 22968 38130
rect 8516 37992 8656 38038
rect 8516 37932 8556 37992
rect 8616 37932 8656 37992
rect 8516 37886 8656 37932
rect 8884 37992 9024 38038
rect 8884 37932 8924 37992
rect 8984 37932 9024 37992
rect 8884 37886 9024 37932
rect 9252 37992 9392 38038
rect 9252 37932 9292 37992
rect 9352 37932 9392 37992
rect 9252 37886 9392 37932
rect 9620 37992 9760 38038
rect 9620 37932 9660 37992
rect 9720 37932 9760 37992
rect 9620 37886 9760 37932
rect 9988 37992 10128 38038
rect 9988 37932 10028 37992
rect 10088 37932 10128 37992
rect 9988 37886 10128 37932
rect 10356 37992 10496 38038
rect 10356 37932 10396 37992
rect 10456 37932 10496 37992
rect 10356 37886 10496 37932
rect 10724 37992 10864 38038
rect 10724 37932 10764 37992
rect 10824 37932 10864 37992
rect 10724 37886 10864 37932
rect 11092 37992 11232 38038
rect 11092 37932 11132 37992
rect 11192 37932 11232 37992
rect 11092 37886 11232 37932
rect 11460 37992 11600 38038
rect 11460 37932 11500 37992
rect 11560 37932 11600 37992
rect 11460 37886 11600 37932
rect 11828 37992 11968 38038
rect 11828 37932 11868 37992
rect 11928 37932 11968 37992
rect 11828 37886 11968 37932
rect 12196 37992 12336 38038
rect 12196 37932 12236 37992
rect 12296 37932 12336 37992
rect 12196 37886 12336 37932
rect 12564 37992 12704 38038
rect 12564 37932 12604 37992
rect 12664 37932 12704 37992
rect 12564 37886 12704 37932
rect 12932 37992 13072 38038
rect 12932 37932 12972 37992
rect 13032 37932 13072 37992
rect 12932 37886 13072 37932
rect 13300 37992 13440 38038
rect 13300 37932 13340 37992
rect 13400 37932 13440 37992
rect 13300 37886 13440 37932
rect 13668 37992 13808 38038
rect 13668 37932 13708 37992
rect 13768 37932 13808 37992
rect 13668 37886 13808 37932
rect 14036 37992 14176 38038
rect 14036 37932 14076 37992
rect 14136 37932 14176 37992
rect 14036 37886 14176 37932
rect 14404 37992 14544 38038
rect 14404 37932 14444 37992
rect 14504 37932 14544 37992
rect 14404 37886 14544 37932
rect 14772 37992 14912 38038
rect 14772 37932 14812 37992
rect 14872 37932 14912 37992
rect 14772 37886 14912 37932
rect 15140 37992 15280 38038
rect 15140 37932 15180 37992
rect 15240 37932 15280 37992
rect 15140 37886 15280 37932
rect 15508 37992 15648 38038
rect 15508 37932 15548 37992
rect 15608 37932 15648 37992
rect 15508 37886 15648 37932
rect 15876 37992 16016 38038
rect 15876 37932 15916 37992
rect 15976 37932 16016 37992
rect 15876 37886 16016 37932
rect 16244 37992 16384 38038
rect 16244 37932 16284 37992
rect 16344 37932 16384 37992
rect 16244 37886 16384 37932
rect 16612 37992 16752 38038
rect 16612 37932 16652 37992
rect 16712 37932 16752 37992
rect 16612 37886 16752 37932
rect 16980 37992 17120 38038
rect 16980 37932 17020 37992
rect 17080 37932 17120 37992
rect 16980 37886 17120 37932
rect 17348 37992 17488 38038
rect 17348 37932 17388 37992
rect 17448 37932 17488 37992
rect 17348 37886 17488 37932
rect 17716 37992 17856 38038
rect 17716 37932 17756 37992
rect 17816 37932 17856 37992
rect 17716 37886 17856 37932
rect 18084 37992 18224 38038
rect 18084 37932 18124 37992
rect 18184 37932 18224 37992
rect 18084 37886 18224 37932
rect 18452 37992 18592 38038
rect 18452 37932 18492 37992
rect 18552 37932 18592 37992
rect 18452 37886 18592 37932
rect 18820 37992 18960 38038
rect 18820 37932 18860 37992
rect 18920 37932 18960 37992
rect 18820 37886 18960 37932
rect 19188 37992 19328 38038
rect 19188 37932 19228 37992
rect 19288 37932 19328 37992
rect 19188 37886 19328 37932
rect 19556 37992 19696 38038
rect 19556 37932 19596 37992
rect 19656 37932 19696 37992
rect 19556 37886 19696 37932
rect 19924 37992 20064 38038
rect 19924 37932 19964 37992
rect 20024 37932 20064 37992
rect 19924 37886 20064 37932
rect 20292 37992 20432 38038
rect 20292 37932 20332 37992
rect 20392 37932 20432 37992
rect 20292 37886 20432 37932
rect 20660 37992 20800 38038
rect 20660 37932 20700 37992
rect 20760 37932 20800 37992
rect 20660 37886 20800 37932
rect 21028 37992 21168 38038
rect 21028 37932 21068 37992
rect 21128 37932 21168 37992
rect 21028 37886 21168 37932
rect 21396 37992 21536 38038
rect 21396 37932 21436 37992
rect 21496 37932 21536 37992
rect 21396 37886 21536 37932
rect 21764 37992 21904 38038
rect 21764 37932 21804 37992
rect 21864 37932 21904 37992
rect 21764 37886 21904 37932
rect 22132 37992 22272 38038
rect 22132 37932 22172 37992
rect 22232 37932 22272 37992
rect 22132 37886 22272 37932
rect 22500 37992 22640 38038
rect 22500 37932 22540 37992
rect 22600 37932 22640 37992
rect 22500 37886 22640 37932
rect 22868 37992 23008 38038
rect 22868 37932 22908 37992
rect 22968 37932 23008 37992
rect 22868 37886 23008 37932
rect 2400 29700 23324 29720
rect 2400 29420 4420 29700
rect 4700 29420 11919 29700
rect 12199 29420 15621 29700
rect 15901 29420 19323 29700
rect 19603 29420 23025 29700
rect 23305 29420 23324 29700
rect 2400 29400 23324 29420
rect 2400 27700 23324 27720
rect 2400 27420 2420 27700
rect 2700 27420 10067 27700
rect 10347 27420 13771 27700
rect 14051 27420 17473 27700
rect 17753 27420 21175 27700
rect 21455 27420 23324 27700
rect 2400 27400 23324 27420
rect 25570 8084 25768 8090
rect 25563 7884 25568 8084
rect 25769 7884 25775 8084
rect 25570 7878 25768 7884
<< via3 >>
rect 788 44962 868 45142
rect 1524 44962 1604 45142
rect 2260 44962 2340 45142
rect 2996 44962 3076 45142
rect 3732 44962 3812 45142
rect 4468 44962 4548 45142
rect 5204 44962 5284 45142
rect 5940 44962 6020 45142
rect 6676 44962 6756 45142
rect 7412 44962 7492 45142
rect 8148 44962 8228 45142
rect 8884 44962 8964 45142
rect 9620 44962 9700 45142
rect 10356 44962 10436 45142
rect 11092 44962 11172 45142
rect 11828 44962 11908 45142
rect 12564 44962 12644 45142
rect 13300 44962 13380 45142
rect 14036 44962 14116 45142
rect 14772 44962 14852 45142
rect 15508 44962 15588 45142
rect 16244 44962 16324 45142
rect 16980 44962 17060 45142
rect 17716 44962 17796 45142
rect 18452 44962 18532 45142
rect 19188 44962 19268 45142
rect 19924 44962 20004 45142
rect 20660 44962 20740 45142
rect 21396 44962 21476 45142
rect 22132 44962 22212 45142
rect 22868 44962 22948 45142
rect 23604 44962 23684 45142
rect 24340 44962 24420 45142
rect 25076 44962 25156 45142
rect 25812 44962 25892 45142
rect 26548 44962 26628 45142
rect 27284 44962 27364 45142
rect 28020 44962 28100 45142
rect 28756 44962 28836 45142
rect 29492 44962 29572 45142
rect 4420 29420 4700 29700
rect 11919 29420 12199 29700
rect 15621 29420 15901 29700
rect 19323 29420 19603 29700
rect 23025 29420 23305 29700
rect 2420 27420 2700 27700
rect 10067 27420 10347 27700
rect 13771 27420 14051 27700
rect 17473 27420 17753 27700
rect 21175 27420 21455 27700
rect 11918 24908 12198 25070
rect 15620 24908 15900 25070
rect 19322 24908 19602 25070
rect 23024 24908 23304 25070
rect 10067 23256 10347 23418
rect 13769 23256 14049 23418
rect 17471 23256 17751 23418
rect 21173 23256 21453 23418
rect 11918 21440 12198 21602
rect 15620 21440 15900 21602
rect 19322 21440 19602 21602
rect 23024 21440 23304 21602
rect 10067 19788 10347 19950
rect 13769 19788 14049 19950
rect 17471 19788 17751 19950
rect 21173 19788 21453 19950
rect 11918 17972 12198 18134
rect 15620 17972 15900 18134
rect 19322 17972 19602 18134
rect 23024 17972 23304 18134
rect 10067 16320 10347 16482
rect 13769 16320 14049 16482
rect 17471 16320 17751 16482
rect 21173 16320 21453 16482
rect 11918 14504 12198 14666
rect 15620 14504 15900 14666
rect 19322 14504 19602 14666
rect 23024 14504 23304 14666
rect 10067 12852 10347 13014
rect 13769 12852 14049 13014
rect 17471 12852 17751 13014
rect 21173 12852 21453 13014
rect 11918 10904 12198 11066
rect 15620 10904 15900 11066
rect 19322 10904 19602 11066
rect 23024 10904 23304 11066
rect 10067 9252 10347 9414
rect 13769 9252 14049 9414
rect 17471 9252 17751 9414
rect 21173 9252 21453 9414
rect 25568 7884 25769 8084
<< metal4 >>
rect 778 45142 878 45152
rect 778 44962 788 45142
rect 868 44962 878 45142
rect 778 44952 878 44962
rect 1514 45142 1614 45152
rect 1514 44962 1524 45142
rect 1604 44962 1614 45142
rect 1514 44952 1614 44962
rect 2250 45142 2350 45152
rect 2250 44962 2260 45142
rect 2340 44962 2350 45142
rect 2250 44952 2350 44962
rect 2986 45142 3086 45152
rect 2986 44962 2996 45142
rect 3076 44962 3086 45142
rect 2986 44952 3086 44962
rect 3722 45142 3822 45152
rect 3722 44962 3732 45142
rect 3812 44962 3822 45142
rect 3722 44952 3822 44962
rect 4458 45142 4558 45152
rect 4458 44962 4468 45142
rect 4548 44962 4558 45142
rect 4458 44952 4558 44962
rect 5194 45142 5294 45152
rect 5194 44962 5204 45142
rect 5284 44962 5294 45142
rect 5194 44952 5294 44962
rect 5930 45142 6030 45152
rect 5930 44962 5940 45142
rect 6020 44962 6030 45142
rect 5930 44952 6030 44962
rect 6666 45142 6766 45152
rect 6666 44962 6676 45142
rect 6756 44962 6766 45142
rect 6666 44952 6766 44962
rect 7402 45142 7502 45152
rect 7402 44962 7412 45142
rect 7492 44962 7502 45142
rect 7402 44952 7502 44962
rect 8138 45142 8238 45152
rect 8138 44962 8148 45142
rect 8228 44962 8238 45142
rect 8138 44952 8238 44962
rect 8874 45142 8974 45152
rect 8874 44962 8884 45142
rect 8964 44962 8974 45142
rect 8874 44952 8974 44962
rect 9610 45142 9710 45152
rect 9610 44962 9620 45142
rect 9700 44962 9710 45142
rect 9610 44952 9710 44962
rect 10346 45142 10446 45152
rect 10346 44962 10356 45142
rect 10436 44962 10446 45142
rect 10346 44952 10446 44962
rect 11082 45142 11182 45152
rect 11082 44962 11092 45142
rect 11172 44962 11182 45142
rect 11082 44952 11182 44962
rect 11818 45142 11918 45152
rect 11818 44962 11828 45142
rect 11908 44962 11918 45142
rect 11818 44952 11918 44962
rect 12554 45142 12654 45152
rect 12554 44962 12564 45142
rect 12644 44962 12654 45142
rect 12554 44952 12654 44962
rect 13290 45142 13390 45152
rect 13290 44962 13300 45142
rect 13380 44962 13390 45142
rect 13290 44952 13390 44962
rect 14026 45142 14126 45152
rect 14026 44962 14036 45142
rect 14116 44962 14126 45142
rect 14026 44952 14126 44962
rect 14762 45142 14862 45152
rect 14762 44962 14772 45142
rect 14852 44962 14862 45142
rect 14762 44952 14862 44962
rect 15498 45142 15598 45152
rect 15498 44962 15508 45142
rect 15588 44962 15598 45142
rect 15498 44952 15598 44962
rect 16234 45142 16334 45152
rect 16234 44962 16244 45142
rect 16324 44962 16334 45142
rect 16234 44952 16334 44962
rect 16970 45142 17070 45152
rect 16970 44962 16980 45142
rect 17060 44962 17070 45142
rect 16970 44952 17070 44962
rect 17706 45142 17806 45152
rect 17706 44962 17716 45142
rect 17796 44962 17806 45142
rect 17706 44952 17806 44962
rect 18442 45142 18542 45152
rect 18442 44962 18452 45142
rect 18532 44962 18542 45142
rect 18442 44952 18542 44962
rect 19178 45142 19278 45152
rect 19178 44962 19188 45142
rect 19268 44962 19278 45142
rect 19178 44952 19278 44962
rect 19914 45142 20014 45152
rect 19914 44962 19924 45142
rect 20004 44962 20014 45142
rect 19914 44952 20014 44962
rect 20650 45142 20750 45152
rect 20650 44962 20660 45142
rect 20740 44962 20750 45142
rect 20650 44952 20750 44962
rect 21386 45142 21486 45152
rect 21386 44962 21396 45142
rect 21476 44962 21486 45142
rect 21386 44952 21486 44962
rect 22122 45142 22222 45152
rect 22122 44962 22132 45142
rect 22212 44962 22222 45142
rect 22122 44952 22222 44962
rect 22858 45142 22958 45152
rect 22858 44962 22868 45142
rect 22948 44962 22958 45142
rect 22858 44952 22958 44962
rect 23594 45142 23694 45152
rect 23594 44962 23604 45142
rect 23684 44962 23694 45142
rect 23594 44952 23694 44962
rect 24330 45142 24430 45152
rect 24330 44962 24340 45142
rect 24420 44962 24430 45142
rect 24330 44952 24430 44962
rect 25066 45142 25166 45152
rect 25066 44962 25076 45142
rect 25156 44962 25166 45142
rect 25066 44952 25166 44962
rect 25802 45142 25902 45152
rect 25802 44962 25812 45142
rect 25892 44962 25902 45142
rect 25802 44952 25902 44962
rect 26538 45142 26638 45152
rect 26538 44962 26548 45142
rect 26628 44962 26638 45142
rect 26538 44952 26638 44962
rect 27274 45142 27374 45152
rect 27274 44962 27284 45142
rect 27364 44962 27374 45142
rect 27274 44952 27374 44962
rect 28010 45142 28110 45152
rect 28010 44962 28020 45142
rect 28100 44962 28110 45142
rect 28010 44952 28110 44962
rect 28746 45142 28846 45152
rect 28746 44962 28756 45142
rect 28836 44962 28846 45142
rect 28746 44952 28846 44962
rect 29482 45142 29582 45152
rect 29482 44962 29492 45142
rect 29572 44962 29582 45142
rect 29482 44952 29582 44962
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 2400 27700 2720 44152
rect 2400 27420 2420 27700
rect 2700 27420 2720 27700
rect 2400 1000 2720 27420
rect 4400 29700 4720 44152
rect 4400 29420 4420 29700
rect 4700 29420 4720 29700
rect 4400 1000 4720 29420
rect 10047 27700 10367 37370
rect 10047 27420 10067 27700
rect 10347 27420 10367 27700
rect 10047 23418 10367 27420
rect 10047 23256 10067 23418
rect 10347 23256 10367 23418
rect 10047 19950 10367 23256
rect 10047 19788 10067 19950
rect 10347 19788 10367 19950
rect 10047 16482 10367 19788
rect 10047 16320 10067 16482
rect 10347 16320 10367 16482
rect 10047 13014 10367 16320
rect 10047 12852 10067 13014
rect 10347 12852 10367 13014
rect 10047 9414 10367 12852
rect 10047 9252 10067 9414
rect 10347 9252 10367 9414
rect 10047 8880 10367 9252
rect 11898 29700 12218 37370
rect 11898 29420 11919 29700
rect 12199 29420 12218 29700
rect 11898 25070 12218 29420
rect 11898 24908 11918 25070
rect 12198 24908 12218 25070
rect 11898 21602 12218 24908
rect 11898 21440 11918 21602
rect 12198 21440 12218 21602
rect 11898 18134 12218 21440
rect 11898 17972 11918 18134
rect 12198 17972 12218 18134
rect 11898 14666 12218 17972
rect 11898 14504 11918 14666
rect 12198 14504 12218 14666
rect 11898 11066 12218 14504
rect 11898 10904 11918 11066
rect 12198 10904 12218 11066
rect 11898 8880 12218 10904
rect 13749 27700 14069 37370
rect 13749 27420 13771 27700
rect 14051 27420 14069 27700
rect 13749 23418 14069 27420
rect 13749 23256 13769 23418
rect 14049 23256 14069 23418
rect 13749 19950 14069 23256
rect 13749 19788 13769 19950
rect 14049 19788 14069 19950
rect 13749 16482 14069 19788
rect 13749 16320 13769 16482
rect 14049 16320 14069 16482
rect 13749 13014 14069 16320
rect 13749 12852 13769 13014
rect 14049 12852 14069 13014
rect 13749 9414 14069 12852
rect 13749 9252 13769 9414
rect 14049 9252 14069 9414
rect 13749 8880 14069 9252
rect 15600 29700 15920 37370
rect 15600 29420 15621 29700
rect 15901 29420 15920 29700
rect 15600 25070 15920 29420
rect 15600 24908 15620 25070
rect 15900 24908 15920 25070
rect 15600 21602 15920 24908
rect 15600 21440 15620 21602
rect 15900 21440 15920 21602
rect 15600 18134 15920 21440
rect 15600 17972 15620 18134
rect 15900 17972 15920 18134
rect 15600 14666 15920 17972
rect 15600 14504 15620 14666
rect 15900 14504 15920 14666
rect 15600 11066 15920 14504
rect 15600 10904 15620 11066
rect 15900 10904 15920 11066
rect 15600 8880 15920 10904
rect 17451 27700 17771 37370
rect 17451 27420 17473 27700
rect 17753 27420 17771 27700
rect 17451 23418 17771 27420
rect 17451 23256 17471 23418
rect 17751 23256 17771 23418
rect 17451 19950 17771 23256
rect 17451 19788 17471 19950
rect 17751 19788 17771 19950
rect 17451 16482 17771 19788
rect 17451 16320 17471 16482
rect 17751 16320 17771 16482
rect 17451 13014 17771 16320
rect 17451 12852 17471 13014
rect 17751 12852 17771 13014
rect 17451 9414 17771 12852
rect 17451 9252 17471 9414
rect 17751 9252 17771 9414
rect 17451 8880 17771 9252
rect 19302 29700 19622 37370
rect 19302 29420 19323 29700
rect 19603 29420 19622 29700
rect 19302 25070 19622 29420
rect 19302 24908 19322 25070
rect 19602 24908 19622 25070
rect 19302 21602 19622 24908
rect 19302 21440 19322 21602
rect 19602 21440 19622 21602
rect 19302 18134 19622 21440
rect 19302 17972 19322 18134
rect 19602 17972 19622 18134
rect 19302 14666 19622 17972
rect 19302 14504 19322 14666
rect 19602 14504 19622 14666
rect 19302 11066 19622 14504
rect 19302 10904 19322 11066
rect 19602 10904 19622 11066
rect 19302 8880 19622 10904
rect 21153 27700 21473 37370
rect 21153 27420 21175 27700
rect 21455 27420 21473 27700
rect 21153 23418 21473 27420
rect 21153 23256 21173 23418
rect 21453 23256 21473 23418
rect 21153 19950 21473 23256
rect 21153 19788 21173 19950
rect 21453 19788 21473 19950
rect 21153 16482 21473 19788
rect 21153 16320 21173 16482
rect 21453 16320 21473 16482
rect 21153 13014 21473 16320
rect 21153 12852 21173 13014
rect 21453 12852 21473 13014
rect 21153 9414 21473 12852
rect 21153 9252 21173 9414
rect 21453 9252 21473 9414
rect 21153 8880 21473 9252
rect 23004 29700 23324 37370
rect 23004 29420 23025 29700
rect 23305 29420 23324 29700
rect 23004 25070 23324 29420
rect 23004 24908 23024 25070
rect 23304 24908 23324 25070
rect 23004 21602 23324 24908
rect 23004 21440 23024 21602
rect 23304 21440 23324 21602
rect 23004 18134 23324 21440
rect 23004 17972 23024 18134
rect 23304 17972 23324 18134
rect 23004 14666 23324 17972
rect 23004 14504 23024 14666
rect 23304 14504 23324 14666
rect 23004 11066 23324 14504
rect 23004 10904 23024 11066
rect 23304 10904 23324 11066
rect 23004 8880 23324 10904
rect 25567 8084 25770 8085
rect 25567 7884 25568 8084
rect 25769 7884 31470 8084
rect 25567 7883 25770 7884
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 200
rect 13648 0 13768 200
rect 18064 0 18184 200
rect 22480 0 22600 200
rect 26896 0 27016 200
rect 31270 0 31470 7884
use encoder  encoder_0
timestamp 1713341310
transform 1 0 7804 0 1 30790
box 514 0 15718 7200
use flash_adc_isolated  flash_adc_isolated_0
timestamp 1713341356
transform -1 0 25768 0 -1 26178
box 0 0 19594 18662
<< labels >>
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal tristate
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal tristate
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal tristate
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal tristate
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal tristate
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal tristate
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal tristate
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal tristate
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal tristate
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal tristate
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal tristate
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal tristate
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal tristate
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal tristate
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal tristate
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal tristate
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal tristate
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal tristate
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal tristate
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal tristate
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal tristate
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal tristate
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal tristate
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal tristate
rlabel metal4 4400 1000 4720 44152 0 VGND
port 52 nsew ground bidirectional
rlabel metal4 2400 1000 2720 44152 0 VPWR
port 51 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
