magic
tech sky130A
magscale 1 2
timestamp 1713023969
<< metal1 >>
rect 1317 6994 1323 7046
rect 1375 7045 1381 7046
rect 5849 7045 5855 7046
rect 1375 6995 5855 7045
rect 1375 6994 1381 6995
rect 5849 6994 5855 6995
rect 5907 6994 5913 7046
rect 10380 6994 10386 7046
rect 10438 7045 10444 7046
rect 14914 7045 14920 7046
rect 10438 6995 14920 7045
rect 10438 6994 10444 6995
rect 14914 6994 14920 6995
rect 14972 6994 14978 7046
rect 5849 -6950 5855 -6898
rect 5907 -6899 5913 -6898
rect 10378 -6899 10384 -6898
rect 5907 -6949 10384 -6899
rect 5907 -6950 5913 -6949
rect 10378 -6950 10384 -6949
rect 10436 -6950 10442 -6898
<< via1 >>
rect 1323 6994 1375 7046
rect 5855 6994 5907 7046
rect 10386 6994 10438 7046
rect 14920 6994 14972 7046
rect 5328 4336 5382 4536
rect 9500 4336 9554 4536
rect 14392 4336 14446 4536
rect 18564 4336 18618 4536
rect 5208 868 5262 1068
rect 9620 868 9674 1068
rect 14272 868 14326 1068
rect 18684 868 18738 1068
rect 5088 -2600 5142 -2400
rect 9740 -2600 9794 -2400
rect 14152 -2600 14206 -2400
rect 18804 -2600 18858 -2400
rect 4968 -6068 5022 -5868
rect 9860 -6068 9914 -5868
rect 14032 -6068 14086 -5868
rect 5855 -6950 5907 -6898
rect 10384 -6950 10436 -6898
<< metal2 >>
rect 5980 10886 6180 10895
rect 1439 10686 1448 10886
rect 1648 10686 1657 10886
rect 858 9536 1058 9545
rect 464 7884 664 7893
rect 464 4286 664 7684
rect 464 820 664 4086
rect 464 -2650 664 620
rect 464 -6118 664 -2850
rect 858 5936 1058 9336
rect 1448 8142 1648 10686
rect 4585 8593 4853 8643
rect 1448 7942 1982 8142
rect 4803 7129 4853 8593
rect 5980 8142 6180 10686
rect 10512 10886 10712 10895
rect 9125 8593 9385 8643
rect 5980 7942 6514 8142
rect 9335 7129 9385 8593
rect 10512 8142 10712 10686
rect 15044 10886 15244 10895
rect 13677 8593 13917 8643
rect 10512 7942 11046 8142
rect 13867 7129 13917 8593
rect 15044 8142 15244 10686
rect 19440 9536 19640 9545
rect 18189 8593 18449 8643
rect 15044 7942 15578 8142
rect 18399 7129 18449 8593
rect 1664 7079 4853 7129
rect 6196 7079 9385 7129
rect 10728 7079 13917 7129
rect 15260 7079 18449 7129
rect 1323 7046 1375 7052
rect 1323 6988 1375 6994
rect 1324 6903 1374 6988
rect 858 2470 1058 5736
rect 1324 3001 1374 4059
rect 858 -1000 1058 2270
rect 1324 -473 1374 593
rect 858 -4473 1058 -1200
rect 1324 -3933 1374 -2869
rect 854 -4663 863 -4473
rect 1053 -4663 1062 -4473
rect 858 -4668 1058 -4663
rect 464 -6327 664 -6318
rect 1249 -6802 1449 -6792
rect 1249 -6982 1259 -6802
rect 1439 -6982 1449 -6802
rect 1664 -6832 1714 7079
rect 5854 7046 5908 7052
rect 5854 6994 5855 7046
rect 5907 6994 5908 7046
rect 5854 6988 5908 6994
rect 5855 6913 5906 6988
rect 5855 6795 5905 6913
rect 5322 4536 5388 4542
rect 5322 4336 5328 4536
rect 5382 4336 5388 4536
rect 5322 4330 5388 4336
rect 5202 1068 5268 1074
rect 5202 868 5208 1068
rect 5262 868 5268 1068
rect 5202 862 5268 868
rect 5082 -2400 5148 -2394
rect 5082 -2600 5088 -2400
rect 5142 -2600 5148 -2400
rect 5082 -2606 5148 -2600
rect 4962 -5868 5028 -5862
rect 4962 -6068 4968 -5868
rect 5022 -6068 5028 -5868
rect 4962 -6074 5028 -6068
rect 4970 -6882 5020 -6074
rect 1249 -6992 1449 -6982
rect 4370 -6932 5020 -6882
rect 4370 -7206 4420 -6932
rect 5090 -6982 5140 -2606
rect 5210 -6739 5260 862
rect 4690 -7032 5140 -6982
rect 5209 -6832 5260 -6739
rect 4690 -7206 4740 -7032
rect 5209 -7082 5259 -6832
rect 5010 -7132 5260 -7082
rect 5010 -7206 5060 -7132
rect 5330 -7206 5380 4330
rect 5856 2997 5906 4063
rect 5856 -465 5906 595
rect 5856 -3937 5906 -2873
rect 5856 -6892 5906 -6771
rect 6196 -6832 6246 7079
rect 10384 7046 10440 7052
rect 10384 6994 10386 7046
rect 10438 6994 10440 7046
rect 10384 6988 10440 6994
rect 10387 6956 10438 6988
rect 10729 6969 10779 7079
rect 14918 7046 14972 7052
rect 14918 6994 14920 7046
rect 14918 6988 14972 6994
rect 10387 6869 10437 6956
rect 10728 6877 10779 6969
rect 14920 6956 14971 6988
rect 14921 6877 14971 6956
rect 9494 4536 9560 4542
rect 9494 4336 9500 4536
rect 9554 4336 9560 4536
rect 9494 4330 9560 4336
rect 9502 -6882 9552 4330
rect 10388 3003 10438 4061
rect 9614 1068 9680 1074
rect 9614 868 9620 1068
rect 9674 868 9680 1068
rect 9614 862 9680 868
rect 5855 -6898 5907 -6892
rect 5855 -6956 5907 -6950
rect 8902 -6932 9552 -6882
rect 8902 -7206 8952 -6932
rect 9622 -6982 9672 862
rect 10388 -469 10438 595
rect 9734 -2400 9800 -2394
rect 9734 -2600 9740 -2400
rect 9794 -2600 9800 -2400
rect 9734 -2606 9800 -2600
rect 9742 -6743 9792 -2606
rect 10388 -3935 10438 -2875
rect 9854 -5868 9920 -5862
rect 9854 -6068 9860 -5868
rect 9914 -6068 9920 -5868
rect 9854 -6074 9920 -6068
rect 9222 -7032 9672 -6982
rect 9741 -6959 9792 -6743
rect 9222 -7206 9272 -7032
rect 9741 -7078 9791 -6959
rect 9741 -7082 9790 -7078
rect 9542 -7132 9790 -7082
rect 9542 -7206 9592 -7132
rect 9862 -7206 9912 -6074
rect 10385 -6892 10435 -6761
rect 10728 -6832 10778 6877
rect 14386 4536 14452 4542
rect 14386 4336 14392 4536
rect 14446 4336 14452 4536
rect 14386 4330 14452 4336
rect 14266 1068 14332 1074
rect 14266 868 14272 1068
rect 14326 868 14332 1068
rect 14266 862 14332 868
rect 14146 -2400 14212 -2394
rect 14146 -2600 14152 -2400
rect 14206 -2600 14212 -2400
rect 14146 -2606 14212 -2600
rect 14026 -5868 14092 -5862
rect 14026 -6068 14032 -5868
rect 14086 -6068 14092 -5868
rect 14026 -6074 14092 -6068
rect 14034 -6882 14084 -6074
rect 10384 -6898 10436 -6892
rect 10384 -6956 10436 -6950
rect 13434 -6932 14084 -6882
rect 4294 -7207 4494 -7206
rect 4294 -7406 4495 -7207
rect 4615 -7406 4816 -7206
rect 4936 -7207 5136 -7206
rect 4935 -7406 5136 -7207
rect 5255 -7406 5456 -7206
rect 8828 -7207 9028 -7206
rect 8827 -7406 9028 -7207
rect 9146 -7406 9347 -7206
rect 9468 -7207 9668 -7206
rect 9467 -7406 9668 -7207
rect 9787 -7406 9988 -7206
rect 13434 -7207 13484 -6932
rect 14154 -6982 14204 -2606
rect 14274 -6844 14324 862
rect 13754 -7032 14204 -6982
rect 14273 -6925 14324 -6844
rect 13754 -7206 13804 -7032
rect 14273 -7082 14323 -6925
rect 14074 -7132 14323 -7082
rect 14074 -7206 14124 -7132
rect 14394 -7206 14444 4330
rect 14920 2997 14970 4061
rect 14920 -467 14970 593
rect 14920 -3448 14970 -3314
rect 15260 -3364 15310 7079
rect 19440 5931 19640 9336
rect 19840 7881 20040 7886
rect 19836 7691 19845 7881
rect 20035 7691 20044 7881
rect 19440 5741 19445 5931
rect 19635 5741 19640 5931
rect 18558 4536 18624 4542
rect 18558 4336 18564 4536
rect 18618 4336 18624 4536
rect 18558 4330 18624 4336
rect 14845 -3458 15045 -3448
rect 14845 -3638 14855 -3458
rect 15035 -3638 15045 -3458
rect 14845 -3648 15045 -3638
rect 18566 -6982 18616 4330
rect 19440 2468 19640 5741
rect 18678 1068 18744 1074
rect 18678 868 18684 1068
rect 18738 868 18744 1068
rect 18678 862 18744 868
rect 18686 -6844 18736 862
rect 19440 -1000 19640 2268
rect 18798 -2400 18864 -2394
rect 18798 -2600 18804 -2400
rect 18858 -2600 18864 -2400
rect 18798 -2606 18864 -2600
rect 18166 -7032 18616 -6982
rect 18685 -6919 18736 -6844
rect 18685 -7014 18735 -6919
rect 18166 -7206 18216 -7032
rect 18685 -7082 18734 -7014
rect 18486 -7132 18734 -7082
rect 13359 -7208 13559 -7207
rect 4295 -7407 4495 -7406
rect 4935 -7407 5135 -7406
rect 8827 -7407 9027 -7406
rect 9467 -7407 9667 -7406
rect 13359 -7407 13560 -7208
rect 13679 -7406 13880 -7206
rect 13998 -7207 14198 -7206
rect 13998 -7406 14199 -7207
rect 14318 -7406 14519 -7206
rect 18091 -7208 18291 -7206
rect 18486 -7207 18536 -7132
rect 18806 -7206 18856 -2606
rect 19440 -4470 19640 -1200
rect 19440 -4679 19640 -4670
rect 19840 4282 20040 7691
rect 19840 818 20040 4082
rect 19840 -2654 20040 618
rect 19840 -6116 20040 -2854
rect 19840 -6325 20040 -6316
rect 18090 -7406 18291 -7208
rect 18411 -7208 18611 -7207
rect 13999 -7407 14199 -7406
rect 13360 -7408 13560 -7407
rect 18090 -7408 18290 -7406
rect 18411 -7407 18612 -7208
rect 18730 -7406 18931 -7206
rect 18412 -7408 18612 -7407
<< via2 >>
rect 1448 10686 1648 10886
rect 5980 10686 6180 10886
rect 858 9336 1058 9536
rect 464 7684 664 7884
rect 464 4086 664 4286
rect 464 620 664 820
rect 464 -2850 664 -2650
rect 10512 10686 10712 10886
rect 15044 10686 15244 10886
rect 19440 9336 19640 9536
rect 858 5736 1058 5936
rect 858 2270 1058 2470
rect 858 -1200 1058 -1000
rect 863 -4663 1053 -4473
rect 464 -6318 664 -6118
rect 1259 -6982 1439 -6802
rect 19845 7691 20035 7881
rect 19445 5741 19635 5931
rect 14855 -3638 15035 -3458
rect 19440 2268 19640 2468
rect 19440 -1200 19640 -1000
rect 19440 -4670 19640 -4470
rect 19840 4082 20040 4282
rect 19840 618 20040 818
rect 19840 -2854 20040 -2654
rect 19840 -6316 20040 -6116
<< metal3 >>
rect 1443 10886 1653 10891
rect 5975 10886 6185 10891
rect 10507 10886 10717 10891
rect 15039 10886 15249 10891
rect 456 10686 1448 10886
rect 1648 10686 5980 10886
rect 6180 10686 10512 10886
rect 10712 10686 15044 10886
rect 15244 10686 20048 10886
rect 1443 10681 1653 10686
rect 5975 10681 6185 10686
rect 10507 10681 10717 10686
rect 15039 10681 15249 10686
rect 853 9538 1063 9541
rect 19435 9538 19645 9541
rect 456 9536 20044 9538
rect 456 9338 858 9536
rect 458 9336 858 9338
rect 1058 9336 19440 9536
rect 19640 9336 20046 9536
rect 853 9331 1063 9336
rect 19435 9331 19645 9336
rect 459 7886 669 7889
rect 458 7884 20046 7886
rect 458 7686 464 7884
rect 459 7684 464 7686
rect 664 7881 20046 7884
rect 664 7691 19845 7881
rect 20035 7691 20046 7881
rect 664 7686 20046 7691
rect 664 7684 669 7686
rect 459 7679 669 7684
rect 853 5938 1063 5941
rect 456 5936 20044 5938
rect 456 5738 858 5936
rect 458 5736 858 5738
rect 1058 5931 20046 5936
rect 1058 5741 19445 5931
rect 19635 5741 20046 5931
rect 1058 5736 20046 5741
rect 853 5731 1063 5736
rect 459 4286 669 4291
rect 19835 4286 20045 4287
rect 458 4086 464 4286
rect 664 4282 20046 4286
rect 664 4086 19840 4282
rect 459 4081 669 4086
rect 19835 4082 19840 4086
rect 20040 4086 20046 4282
rect 20040 4082 20045 4086
rect 19835 4077 20045 4082
rect 853 2470 1063 2475
rect 19435 2470 19645 2473
rect 456 2270 858 2470
rect 1058 2468 20044 2470
rect 1058 2270 19440 2468
rect 458 2268 19440 2270
rect 19640 2268 20046 2468
rect 853 2265 1063 2268
rect 19435 2263 19645 2268
rect 459 820 669 825
rect 459 818 464 820
rect 458 620 464 818
rect 664 818 669 820
rect 19835 818 20045 823
rect 664 620 19840 818
rect 458 618 19840 620
rect 20040 618 20046 818
rect 459 615 669 618
rect 19835 613 20045 618
rect 853 -998 1063 -995
rect 19435 -998 19645 -995
rect 456 -1000 20044 -998
rect 456 -1198 858 -1000
rect 458 -1200 858 -1198
rect 1058 -1200 19440 -1000
rect 19640 -1200 20046 -1000
rect 853 -1205 1063 -1200
rect 19435 -1205 19645 -1200
rect 459 -2650 669 -2645
rect 19835 -2650 20045 -2649
rect 458 -2850 464 -2650
rect 664 -2654 20046 -2650
rect 664 -2850 19840 -2654
rect 459 -2855 669 -2850
rect 19835 -2854 19840 -2850
rect 20040 -2850 20046 -2654
rect 20040 -2854 20045 -2850
rect 19835 -2859 20045 -2854
rect 14845 -3458 15045 -3448
rect 14845 -3638 14855 -3458
rect 15035 -3638 15045 -3458
rect 14845 -4466 15045 -3638
rect 19435 -4466 19645 -4465
rect 456 -4468 20044 -4466
rect 456 -4470 20046 -4468
rect 456 -4473 19440 -4470
rect 456 -4663 863 -4473
rect 1053 -4663 19440 -4473
rect 456 -4666 19440 -4663
rect 458 -4668 19440 -4666
rect 19435 -4670 19440 -4668
rect 19640 -4668 20046 -4470
rect 19640 -4670 19645 -4668
rect 19435 -4675 19645 -4670
rect 459 -6118 669 -6113
rect 19835 -6116 20045 -6111
rect 19835 -6118 19840 -6116
rect 458 -6318 464 -6118
rect 664 -6316 19840 -6118
rect 20040 -6118 20045 -6116
rect 20040 -6316 20046 -6118
rect 664 -6318 20046 -6316
rect 459 -6323 669 -6318
rect 1249 -6802 1449 -6318
rect 19835 -6321 20045 -6318
rect 1249 -6982 1259 -6802
rect 1439 -6982 1449 -6802
rect 1249 -6992 1449 -6982
use ladder_rung  ladder_rung_0
timestamp 1713023969
transform 1 0 56 0 1 -4974
box 1092 -1858 5604 1538
use ladder_rung  ladder_rung_1
timestamp 1713023969
transform 1 0 56 0 1 -1506
box 1092 -1858 5604 1538
use ladder_rung  ladder_rung_2
timestamp 1713023969
transform 1 0 56 0 1 1962
box 1092 -1858 5604 1538
use ladder_rung  ladder_rung_3
timestamp 1713023969
transform 1 0 56 0 1 5430
box 1092 -1858 5604 1538
use ladder_rung  ladder_rung_4
timestamp 1713023969
transform 1 0 4588 0 1 5430
box 1092 -1858 5604 1538
use ladder_rung  ladder_rung_5
timestamp 1713023969
transform 1 0 4588 0 1 1962
box 1092 -1858 5604 1538
use ladder_rung  ladder_rung_6
timestamp 1713023969
transform 1 0 4588 0 1 -1506
box 1092 -1858 5604 1538
use ladder_rung  ladder_rung_7
timestamp 1713023969
transform 1 0 4588 0 1 -4974
box 1092 -1858 5604 1538
use ladder_rung  ladder_rung_8
timestamp 1713023969
transform 1 0 9120 0 1 -4974
box 1092 -1858 5604 1538
use ladder_rung  ladder_rung_9
timestamp 1713023969
transform 1 0 9120 0 1 -1506
box 1092 -1858 5604 1538
use ladder_rung  ladder_rung_10
timestamp 1713023969
transform 1 0 9120 0 1 1962
box 1092 -1858 5604 1538
use ladder_rung  ladder_rung_11
timestamp 1713023969
transform 1 0 9120 0 1 5430
box 1092 -1858 5604 1538
use ladder_rung  ladder_rung_12
timestamp 1713023969
transform 1 0 13652 0 1 5430
box 1092 -1858 5604 1538
use ladder_rung  ladder_rung_13
timestamp 1713023969
transform 1 0 13652 0 1 1962
box 1092 -1858 5604 1538
use ladder_rung  ladder_rung_14
timestamp 1713023969
transform 1 0 13652 0 1 -1506
box 1092 -1858 5604 1538
use vfollower  vfollower_0
timestamp 1713023969
transform 1 0 1414 0 1 8370
box 368 -1198 3296 2198
use vfollower  vfollower_1
timestamp 1713023969
transform 1 0 5946 0 1 8370
box 368 -1198 3296 2198
use vfollower  vfollower_2
timestamp 1713023969
transform 1 0 10478 0 1 8370
box 368 -1198 3296 2198
use vfollower  vfollower_3
timestamp 1713023969
transform 1 0 15010 0 1 8370
box 368 -1198 3296 2198
<< labels >>
flabel metal2 4294 -7406 4494 -7206 0 FreeSans 256 0 0 0 OUT0
port 16 nsew
flabel metal2 4616 -7406 4816 -7206 0 FreeSans 256 0 0 0 OUT1
port 15 nsew
flabel metal2 4936 -7406 5136 -7206 0 FreeSans 256 0 0 0 OUT2
port 14 nsew
flabel metal2 5256 -7406 5456 -7206 0 FreeSans 256 0 0 0 OUT3
port 13 nsew
flabel metal2 8828 -7406 9028 -7206 0 FreeSans 256 0 0 0 OUT4
port 12 nsew
flabel metal2 9146 -7406 9346 -7206 0 FreeSans 256 0 0 0 OUT5
port 11 nsew
flabel metal2 9468 -7406 9668 -7206 0 FreeSans 256 0 0 0 OUT6
port 10 nsew
flabel metal2 9788 -7406 9988 -7206 0 FreeSans 256 0 0 0 OUT7
port 9 nsew
flabel metal2 13360 -7408 13560 -7208 0 FreeSans 256 0 0 0 OUT8
port 8 nsew
flabel metal2 13680 -7406 13880 -7206 0 FreeSans 256 0 0 0 OUT9
port 7 nsew
flabel metal2 13998 -7406 14198 -7206 0 FreeSans 256 0 0 0 OUT10
port 6 nsew
flabel metal2 14318 -7406 14518 -7206 0 FreeSans 256 0 0 0 OUT11
port 5 nsew
flabel metal2 18090 -7408 18290 -7208 0 FreeSans 256 0 0 0 OUT12
port 4 nsew
flabel metal2 18412 -7408 18612 -7208 0 FreeSans 256 0 0 0 OUT13
port 3 nsew
flabel metal2 18730 -7406 18930 -7206 0 FreeSans 256 0 0 0 OUT14
port 2 nsew
flabel metal3 458 7686 20046 7886 0 FreeSans 256 0 0 0 VSS
port 17 nsew
flabel metal3 456 9338 20044 9538 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal3 456 5738 20044 5938 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal3 458 4086 20046 4286 0 FreeSans 256 0 0 0 VSS
port 17 nsew
flabel metal3 456 2270 20044 2470 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal3 458 618 20046 818 0 FreeSans 256 0 0 0 VSS
port 17 nsew
flabel metal3 458 -2850 20046 -2650 0 FreeSans 256 0 0 0 VSS
port 17 nsew
flabel metal3 456 -1198 20044 -998 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal3 458 -6318 20046 -6118 0 FreeSans 256 0 0 0 VSS
port 17 nsew
flabel metal3 456 -4666 20044 -4466 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal3 456 10686 20048 10886 0 FreeSans 256 0 0 0 IN
port 1 nsew
<< end >>
