magic
tech sky130A
magscale 1 2
timestamp 1712769939
<< dnwell >>
rect 440 300 19376 18582
<< nwell >>
rect 360 18376 19456 18662
rect 360 506 646 18376
rect 19170 506 19456 18376
rect 360 220 19456 506
<< nsubdiff >>
rect 397 18605 19419 18625
rect 397 18571 477 18605
rect 19339 18571 19419 18605
rect 397 18551 19419 18571
rect 397 18545 471 18551
rect 397 337 417 18545
rect 451 337 471 18545
rect 397 331 471 337
rect 19345 18545 19419 18551
rect 19345 337 19365 18545
rect 19399 337 19419 18545
rect 19345 331 19419 337
rect 397 311 19419 331
rect 397 277 477 311
rect 19339 277 19419 311
rect 397 257 19419 277
<< nsubdiffcont >>
rect 477 18571 19339 18605
rect 417 337 451 18545
rect 19365 337 19399 18545
rect 477 277 19339 311
<< locali >>
rect 417 18571 477 18605
rect 19339 18571 19399 18605
rect 417 18545 451 18571
rect 417 311 451 337
rect 19365 18545 19399 18571
rect 19365 311 19399 337
rect 417 277 477 311
rect 19339 277 19399 311
<< metal2 >>
rect 8 11694 208 15092
rect 8 8228 208 11494
rect 8 4758 208 8028
rect 8 1290 208 4558
rect 402 13344 602 16744
rect 18984 13339 19184 16744
rect 402 9878 602 13144
rect 402 6408 602 9678
rect 402 2935 602 6208
rect 18984 9876 19184 13149
rect 18984 6408 19184 9676
rect 18984 2938 19184 6208
rect 19384 11690 19584 15099
rect 19384 8226 19584 11490
rect 19384 4754 19584 8026
rect 19384 1292 19584 4554
rect 3838 2 4038 202
rect 4159 2 4360 202
rect 4480 2 4680 202
rect 4799 2 5000 202
rect 8371 1 8571 201
rect 8690 2 8891 202
rect 9012 2 9212 202
rect 9331 2 9532 202
rect 12903 1 13103 201
rect 13223 2 13424 202
rect 13542 2 13742 202
rect 13862 2 14063 202
rect 17635 2 17835 202
rect 17955 1 18155 201
rect 18274 2 18475 202
<< via2 >>
rect 402 16744 602 16944
rect 8 15092 208 15292
rect 8 11494 208 11694
rect 8 8028 208 8228
rect 8 4558 208 4758
rect 402 13144 602 13344
rect 18984 16744 19184 16944
rect 19389 15099 19579 15289
rect 18989 13149 19179 13339
rect 402 9678 602 9878
rect 402 6208 602 6408
rect 18984 9676 19184 9876
rect 18984 6208 19184 6408
rect 407 2745 597 2935
rect 18984 2738 19184 2938
rect 19384 11490 19584 11690
rect 19384 8026 19584 8226
rect 19384 4554 19584 4754
rect 19384 1092 19584 1292
<< metal3 >>
rect 0 18094 19592 18294
rect 0 16944 19592 16946
rect 0 16746 402 16944
rect 602 16746 18984 16944
rect 19184 16746 19592 16944
rect 2 15292 19594 15294
rect 2 15094 8 15292
rect 208 15289 19594 15292
rect 208 15099 19389 15289
rect 19579 15099 19594 15289
rect 208 15094 19594 15099
rect 0 13344 19592 13346
rect 0 13146 402 13344
rect 602 13339 19592 13344
rect 602 13149 18989 13339
rect 19179 13149 19592 13339
rect 602 13146 19592 13149
rect 2 11494 8 11694
rect 208 11690 19594 11694
rect 208 11494 19384 11690
rect 19584 11494 19594 11690
rect 0 9678 402 9878
rect 602 9876 19592 9878
rect 602 9678 18984 9876
rect 19184 9678 19592 9876
rect 2 8028 8 8226
rect 208 8028 19384 8226
rect 2 8026 19384 8028
rect 19584 8026 19594 8226
rect 0 6408 19592 6410
rect 0 6210 402 6408
rect 602 6210 18984 6408
rect 19184 6210 19592 6408
rect 2 4558 8 4758
rect 208 4754 19594 4758
rect 208 4558 19384 4754
rect 19584 4558 19594 4754
rect 0 2938 19592 2942
rect 0 2935 18984 2938
rect 0 2745 407 2935
rect 597 2745 18984 2935
rect 0 2742 18984 2745
rect 19184 2742 19592 2938
rect 3 1290 213 1295
rect 2 1092 19384 1290
rect 19584 1092 19594 1290
rect 2 1090 19594 1092
rect 3 1085 213 1090
use flash_adc  flash_adc_0
timestamp 1712769939
transform 1 0 -456 0 1 7408
box 456 -7408 20048 10895
<< labels >>
flabel metal2 3838 2 4038 202 0 FreeSans 256 0 0 0 OUT0
port 16 nsew
flabel metal2 4160 2 4360 202 0 FreeSans 256 0 0 0 OUT1
port 15 nsew
flabel metal2 4480 2 4680 202 0 FreeSans 256 0 0 0 OUT2
port 14 nsew
flabel metal2 4800 2 5000 202 0 FreeSans 256 0 0 0 OUT3
port 13 nsew
flabel metal2 8372 2 8572 202 0 FreeSans 256 0 0 0 OUT4
port 12 nsew
flabel metal2 8690 2 8890 202 0 FreeSans 256 0 0 0 OUT5
port 11 nsew
flabel metal2 9012 2 9212 202 0 FreeSans 256 0 0 0 OUT6
port 10 nsew
flabel metal2 9332 2 9532 202 0 FreeSans 256 0 0 0 OUT7
port 9 nsew
flabel metal2 12904 0 13104 200 0 FreeSans 256 0 0 0 OUT8
port 8 nsew
flabel metal2 13224 2 13424 202 0 FreeSans 256 0 0 0 OUT9
port 7 nsew
flabel metal2 13542 2 13742 202 0 FreeSans 256 0 0 0 OUT10
port 6 nsew
flabel metal2 13862 2 14062 202 0 FreeSans 256 0 0 0 OUT11
port 5 nsew
flabel metal2 17634 0 17834 200 0 FreeSans 256 0 0 0 OUT12
port 4 nsew
flabel metal2 17956 0 18156 200 0 FreeSans 256 0 0 0 OUT13
port 3 nsew
flabel metal2 18274 2 18474 202 0 FreeSans 256 0 0 0 OUT14
port 2 nsew
flabel metal3 2 15094 19590 15294 0 FreeSans 256 0 0 0 VSS
port 17 nsew
flabel metal3 0 16746 19588 16946 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal3 0 13146 19588 13346 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal3 2 11494 19590 11694 0 FreeSans 256 0 0 0 VSS
port 17 nsew
flabel metal3 0 9678 19588 9878 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal3 2 8026 19590 8226 0 FreeSans 256 0 0 0 VSS
port 17 nsew
flabel metal3 2 4558 19590 4758 0 FreeSans 256 0 0 0 VSS
port 17 nsew
flabel metal3 0 6210 19588 6410 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal3 2 1090 19590 1290 0 FreeSans 256 0 0 0 VSS
port 17 nsew
flabel metal3 0 2742 19588 2942 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal3 0 18094 19592 18294 0 FreeSans 256 0 0 0 IN
port 1 nsew
<< end >>
