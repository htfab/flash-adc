magic
tech sky130A
magscale 1 2
timestamp 1712769939
<< viali >>
rect 1409 6409 1443 6443
rect 1961 6409 1995 6443
rect 2421 6409 2455 6443
rect 2789 6409 2823 6443
rect 3341 6409 3375 6443
rect 3893 6409 3927 6443
rect 4537 6409 4571 6443
rect 5181 6409 5215 6443
rect 5917 6409 5951 6443
rect 6377 6409 6411 6443
rect 6653 6409 6687 6443
rect 7205 6409 7239 6443
rect 7665 6409 7699 6443
rect 9229 6409 9263 6443
rect 12081 6409 12115 6443
rect 4261 6341 4295 6375
rect 5549 6341 5583 6375
rect 9689 6341 9723 6375
rect 13829 6341 13863 6375
rect 8769 6273 8803 6307
rect 11069 6273 11103 6307
rect 12633 6273 12667 6307
rect 14657 6273 14691 6307
rect 1133 6205 1167 6239
rect 1777 6205 1811 6239
rect 2237 6205 2271 6239
rect 2605 6205 2639 6239
rect 3525 6205 3559 6239
rect 3709 6205 3743 6239
rect 4077 6205 4111 6239
rect 4721 6205 4755 6239
rect 5365 6205 5399 6239
rect 6101 6205 6135 6239
rect 6193 6205 6227 6239
rect 6837 6205 6871 6239
rect 7389 6205 7423 6239
rect 7849 6205 7883 6239
rect 9045 6205 9079 6239
rect 9873 6205 9907 6239
rect 10241 6205 10275 6239
rect 10609 6205 10643 6239
rect 11621 6205 11655 6239
rect 14013 6205 14047 6239
rect 4905 6137 4939 6171
rect 9505 6137 9539 6171
rect 12357 6137 12391 6171
rect 14565 6137 14599 6171
rect 10057 6069 10091 6103
rect 10425 6069 10459 6103
rect 12817 6069 12851 6103
rect 12909 6069 12943 6103
rect 13277 6069 13311 6103
rect 14105 6069 14139 6103
rect 14473 6069 14507 6103
rect 1133 5865 1167 5899
rect 1593 5865 1627 5899
rect 3985 5865 4019 5899
rect 5641 5865 5675 5899
rect 6745 5865 6779 5899
rect 7113 5865 7147 5899
rect 9045 5865 9079 5899
rect 10977 5865 11011 5899
rect 11805 5865 11839 5899
rect 12173 5865 12207 5899
rect 3249 5797 3283 5831
rect 6285 5797 6319 5831
rect 10149 5797 10183 5831
rect 12817 5797 12851 5831
rect 1317 5729 1351 5763
rect 1409 5729 1443 5763
rect 3525 5729 3559 5763
rect 5273 5729 5307 5763
rect 6377 5729 6411 5763
rect 7205 5729 7239 5763
rect 8217 5729 8251 5763
rect 8953 5729 8987 5763
rect 10793 5729 10827 5763
rect 11345 5729 11379 5763
rect 11437 5729 11471 5763
rect 13369 5729 13403 5763
rect 13921 5729 13955 5763
rect 14381 5729 14415 5763
rect 3801 5661 3835 5695
rect 5089 5661 5123 5695
rect 5181 5661 5215 5695
rect 6101 5661 6135 5695
rect 7021 5661 7055 5695
rect 8493 5661 8527 5695
rect 9229 5661 9263 5695
rect 10241 5661 10275 5695
rect 10333 5661 10367 5695
rect 11529 5661 11563 5695
rect 12265 5661 12299 5695
rect 12357 5661 12391 5695
rect 14013 5661 14047 5695
rect 14105 5661 14139 5695
rect 14565 5661 14599 5695
rect 2881 5593 2915 5627
rect 3433 5593 3467 5627
rect 3617 5593 3651 5627
rect 8585 5593 8619 5627
rect 9781 5593 9815 5627
rect 3249 5525 3283 5559
rect 7573 5525 7607 5559
rect 10609 5525 10643 5559
rect 13553 5525 13587 5559
rect 4813 5321 4847 5355
rect 10977 5321 11011 5355
rect 11345 5321 11379 5355
rect 12265 5321 12299 5355
rect 11621 5253 11655 5287
rect 5457 5185 5491 5219
rect 10149 5185 10183 5219
rect 12817 5185 12851 5219
rect 14013 5185 14047 5219
rect 14289 5185 14323 5219
rect 2329 5117 2363 5151
rect 2605 5117 2639 5151
rect 2789 5117 2823 5151
rect 2973 5117 3007 5151
rect 3065 5117 3099 5151
rect 5181 5117 5215 5151
rect 6009 5117 6043 5151
rect 6745 5117 6779 5151
rect 7389 5117 7423 5151
rect 10793 5117 10827 5151
rect 11529 5117 11563 5151
rect 11805 5117 11839 5151
rect 12081 5117 12115 5151
rect 13277 5117 13311 5151
rect 13645 5117 13679 5151
rect 7205 5049 7239 5083
rect 10241 5049 10275 5083
rect 12633 5049 12667 5083
rect 2145 4981 2179 5015
rect 5273 4981 5307 5015
rect 5825 4981 5859 5015
rect 6653 4981 6687 5015
rect 10333 4981 10367 5015
rect 10701 4981 10735 5015
rect 11897 4981 11931 5015
rect 12725 4981 12759 5015
rect 13093 4981 13127 5015
rect 13737 4981 13771 5015
rect 3893 4777 3927 4811
rect 4261 4777 4295 4811
rect 4905 4777 4939 4811
rect 7389 4777 7423 4811
rect 7849 4777 7883 4811
rect 10977 4777 11011 4811
rect 13829 4777 13863 4811
rect 8217 4709 8251 4743
rect 13277 4709 13311 4743
rect 2329 4641 2363 4675
rect 4813 4641 4847 4675
rect 6009 4641 6043 4675
rect 6193 4641 6227 4675
rect 7757 4641 7791 4675
rect 9020 4641 9054 4675
rect 9137 4641 9171 4675
rect 9873 4641 9907 4675
rect 10149 4641 10183 4675
rect 10333 4641 10367 4675
rect 11345 4641 11379 4675
rect 11897 4641 11931 4675
rect 13185 4641 13219 4675
rect 14013 4641 14047 4675
rect 14933 4641 14967 4675
rect 2513 4573 2547 4607
rect 2605 4573 2639 4607
rect 4353 4573 4387 4607
rect 4445 4573 4479 4607
rect 5825 4573 5859 4607
rect 7941 4573 7975 4607
rect 8861 4573 8895 4607
rect 9413 4573 9447 4607
rect 10057 4573 10091 4607
rect 10517 4573 10551 4607
rect 11437 4573 11471 4607
rect 11621 4573 11655 4607
rect 12449 4573 12483 4607
rect 13369 4573 13403 4607
rect 14473 4573 14507 4607
rect 2145 4505 2179 4539
rect 12817 4437 12851 4471
rect 3709 4233 3743 4267
rect 10609 4233 10643 4267
rect 11713 4233 11747 4267
rect 2513 4165 2547 4199
rect 6929 4165 6963 4199
rect 9137 4165 9171 4199
rect 2237 4097 2271 4131
rect 3341 4097 3375 4131
rect 4261 4097 4295 4131
rect 4721 4097 4755 4131
rect 6009 4097 6043 4131
rect 6423 4097 6457 4131
rect 7322 4097 7356 4131
rect 8585 4097 8619 4131
rect 8677 4097 8711 4131
rect 10057 4097 10091 4131
rect 10885 4097 10919 4131
rect 12357 4097 12391 4131
rect 13001 4097 13035 4131
rect 13093 4097 13127 4131
rect 14105 4097 14139 4131
rect 14749 4097 14783 4131
rect 2145 4029 2179 4063
rect 3433 4029 3467 4063
rect 4077 4029 4111 4063
rect 6285 4029 6319 4063
rect 7205 4029 7239 4063
rect 7481 4029 7515 4063
rect 8125 4029 8159 4063
rect 9413 4029 9447 4063
rect 10149 4029 10183 4063
rect 10241 4029 10275 4063
rect 12909 4029 12943 4063
rect 13921 4029 13955 4063
rect 15025 4029 15059 4063
rect 4997 3961 5031 3995
rect 8769 3961 8803 3995
rect 12081 3961 12115 3995
rect 3893 3893 3927 3927
rect 4905 3893 4939 3927
rect 5365 3893 5399 3927
rect 5457 3893 5491 3927
rect 5825 3893 5859 3927
rect 5917 3893 5951 3927
rect 9229 3893 9263 3927
rect 10977 3893 11011 3927
rect 11069 3893 11103 3927
rect 11437 3893 11471 3927
rect 12173 3893 12207 3927
rect 12541 3893 12575 3927
rect 13553 3893 13587 3927
rect 14013 3893 14047 3927
rect 3433 3689 3467 3723
rect 8861 3689 8895 3723
rect 10241 3689 10275 3723
rect 15025 3689 15059 3723
rect 12541 3621 12575 3655
rect 3801 3553 3835 3587
rect 4997 3553 5031 3587
rect 5181 3553 5215 3587
rect 5825 3553 5859 3587
rect 8769 3553 8803 3587
rect 9597 3553 9631 3587
rect 9781 3553 9815 3587
rect 11805 3553 11839 3587
rect 11989 3553 12023 3587
rect 13185 3553 13219 3587
rect 13369 3553 13403 3587
rect 14105 3553 14139 3587
rect 3893 3485 3927 3519
rect 4077 3485 4111 3519
rect 9045 3485 9079 3519
rect 14222 3485 14256 3519
rect 14381 3485 14415 3519
rect 5365 3417 5399 3451
rect 13829 3417 13863 3451
rect 4813 3349 4847 3383
rect 6009 3349 6043 3383
rect 8401 3349 8435 3383
rect 9873 3349 9907 3383
rect 12081 3349 12115 3383
rect 4997 3145 5031 3179
rect 6377 3145 6411 3179
rect 10425 3145 10459 3179
rect 11345 3145 11379 3179
rect 13553 3145 13587 3179
rect 13369 3077 13403 3111
rect 14381 3077 14415 3111
rect 14657 3077 14691 3111
rect 4353 3009 4387 3043
rect 7113 3009 7147 3043
rect 9229 3009 9263 3043
rect 9622 3009 9656 3043
rect 10793 3009 10827 3043
rect 11713 3009 11747 3043
rect 12173 3009 12207 3043
rect 12449 3009 12483 3043
rect 14105 3009 14139 3043
rect 5825 2941 5859 2975
rect 5917 2941 5951 2975
rect 6101 2941 6135 2975
rect 6929 2941 6963 2975
rect 7021 2941 7055 2975
rect 8585 2941 8619 2975
rect 8769 2941 8803 2975
rect 9505 2941 9539 2975
rect 9781 2941 9815 2975
rect 10885 2941 10919 2975
rect 11069 2941 11103 2975
rect 11529 2941 11563 2975
rect 12566 2941 12600 2975
rect 12725 2941 12759 2975
rect 14013 2941 14047 2975
rect 14565 2941 14599 2975
rect 14841 2941 14875 2975
rect 4537 2805 4571 2839
rect 4629 2805 4663 2839
rect 6561 2805 6595 2839
rect 13921 2805 13955 2839
rect 2329 2601 2363 2635
rect 6469 2601 6503 2635
rect 11621 2601 11655 2635
rect 13185 2601 13219 2635
rect 6561 2533 6595 2567
rect 7573 2533 7607 2567
rect 8309 2533 8343 2567
rect 14565 2533 14599 2567
rect 3132 2465 3166 2499
rect 3249 2465 3283 2499
rect 4031 2465 4065 2499
rect 7389 2465 7423 2499
rect 8125 2465 8159 2499
rect 10701 2465 10735 2499
rect 11161 2465 11195 2499
rect 11345 2465 11379 2499
rect 13645 2465 13679 2499
rect 14657 2465 14691 2499
rect 2973 2397 3007 2431
rect 4169 2397 4203 2431
rect 7757 2397 7791 2431
rect 11069 2397 11103 2431
rect 13829 2397 13863 2431
rect 14749 2397 14783 2431
rect 3525 2329 3559 2363
rect 7205 2329 7239 2363
rect 10517 2329 10551 2363
rect 13553 2261 13587 2295
rect 14197 2261 14231 2295
rect 4445 2057 4479 2091
rect 9045 2057 9079 2091
rect 10977 2057 11011 2091
rect 12817 2057 12851 2091
rect 14657 2057 14691 2091
rect 5641 1989 5675 2023
rect 14105 1989 14139 2023
rect 3525 1921 3559 1955
rect 5089 1921 5123 1955
rect 6101 1921 6135 1955
rect 9965 1921 9999 1955
rect 11529 1921 11563 1955
rect 12357 1921 12391 1955
rect 3617 1853 3651 1887
rect 5248 1853 5282 1887
rect 5365 1853 5399 1887
rect 6285 1853 6319 1887
rect 8493 1853 8527 1887
rect 8585 1853 8619 1887
rect 8769 1853 8803 1887
rect 9781 1853 9815 1887
rect 9873 1853 9907 1887
rect 11437 1853 11471 1887
rect 14289 1853 14323 1887
rect 14565 1853 14599 1887
rect 14841 1853 14875 1887
rect 8125 1785 8159 1819
rect 12173 1785 12207 1819
rect 12725 1785 12759 1819
rect 3249 1717 3283 1751
rect 8033 1717 8067 1751
rect 9413 1717 9447 1751
rect 11345 1717 11379 1751
rect 11805 1717 11839 1751
rect 12265 1717 12299 1751
rect 14381 1717 14415 1751
rect 3801 1513 3835 1547
rect 6193 1513 6227 1547
rect 7021 1513 7055 1547
rect 7389 1513 7423 1547
rect 12541 1513 12575 1547
rect 13369 1513 13403 1547
rect 14381 1513 14415 1547
rect 14657 1513 14691 1547
rect 11529 1445 11563 1479
rect 13001 1445 13035 1479
rect 13553 1445 13587 1479
rect 2789 1377 2823 1411
rect 3433 1377 3467 1411
rect 4629 1377 4663 1411
rect 5273 1377 5307 1411
rect 6561 1377 6595 1411
rect 8217 1377 8251 1411
rect 10517 1377 10551 1411
rect 12909 1377 12943 1411
rect 14565 1377 14599 1411
rect 14841 1377 14875 1411
rect 2881 1309 2915 1343
rect 3157 1309 3191 1343
rect 3341 1309 3375 1343
rect 4721 1309 4755 1343
rect 5365 1309 5399 1343
rect 6653 1309 6687 1343
rect 6837 1309 6871 1343
rect 7481 1309 7515 1343
rect 7573 1309 7607 1343
rect 8125 1309 8159 1343
rect 10609 1309 10643 1343
rect 13093 1309 13127 1343
rect 13737 1309 13771 1343
rect 4997 1241 5031 1275
rect 11345 1241 11379 1275
rect 13921 1241 13955 1275
rect 5641 1173 5675 1207
rect 8493 1173 8527 1207
rect 10149 1173 10183 1207
rect 1133 969 1167 1003
rect 3433 969 3467 1003
rect 4169 969 4203 1003
rect 5181 969 5215 1003
rect 6285 969 6319 1003
rect 7205 969 7239 1003
rect 8033 969 8067 1003
rect 9689 969 9723 1003
rect 10241 969 10275 1003
rect 11253 969 11287 1003
rect 12265 969 12299 1003
rect 13277 969 13311 1003
rect 14197 969 14231 1003
rect 14841 969 14875 1003
rect 2145 901 2179 935
rect 5917 833 5951 867
rect 9137 833 9171 867
rect 14105 833 14139 867
rect 949 765 983 799
rect 1961 765 1995 799
rect 3249 765 3283 799
rect 3985 765 4019 799
rect 4997 765 5031 799
rect 6009 765 6043 799
rect 6469 765 6503 799
rect 7021 765 7055 799
rect 8217 765 8251 799
rect 9229 765 9263 799
rect 9505 765 9539 799
rect 10057 765 10091 799
rect 11069 765 11103 799
rect 12081 765 12115 799
rect 13093 765 13127 799
rect 13737 765 13771 799
rect 13921 765 13955 799
rect 14381 765 14415 799
rect 15025 765 15059 799
rect 6653 629 6687 663
rect 8861 629 8895 663
rect 14565 629 14599 663
<< metal1 >>
rect 7466 6740 7472 6792
rect 7524 6780 7530 6792
rect 10870 6780 10876 6792
rect 7524 6752 10876 6780
rect 7524 6740 7530 6752
rect 10870 6740 10876 6752
rect 10928 6740 10934 6792
rect 12250 6740 12256 6792
rect 12308 6780 12314 6792
rect 15010 6780 15016 6792
rect 12308 6752 15016 6780
rect 12308 6740 12314 6752
rect 15010 6740 15016 6752
rect 15068 6740 15074 6792
rect 7098 6672 7104 6724
rect 7156 6712 7162 6724
rect 15654 6712 15660 6724
rect 7156 6684 15660 6712
rect 7156 6672 7162 6684
rect 15654 6672 15660 6684
rect 15712 6672 15718 6724
rect 8110 6604 8116 6656
rect 8168 6644 8174 6656
rect 11974 6644 11980 6656
rect 8168 6616 11980 6644
rect 8168 6604 8174 6616
rect 11974 6604 11980 6616
rect 12032 6604 12038 6656
rect 12894 6604 12900 6656
rect 12952 6644 12958 6656
rect 15562 6644 15568 6656
rect 12952 6616 15568 6644
rect 12952 6604 12958 6616
rect 15562 6604 15568 6616
rect 15620 6604 15626 6656
rect 552 6554 15364 6576
rect 552 6502 2249 6554
rect 2301 6502 2313 6554
rect 2365 6502 2377 6554
rect 2429 6502 2441 6554
rect 2493 6502 2505 6554
rect 2557 6502 5951 6554
rect 6003 6502 6015 6554
rect 6067 6502 6079 6554
rect 6131 6502 6143 6554
rect 6195 6502 6207 6554
rect 6259 6502 9653 6554
rect 9705 6502 9717 6554
rect 9769 6502 9781 6554
rect 9833 6502 9845 6554
rect 9897 6502 9909 6554
rect 9961 6502 13355 6554
rect 13407 6502 13419 6554
rect 13471 6502 13483 6554
rect 13535 6502 13547 6554
rect 13599 6502 13611 6554
rect 13663 6502 15364 6554
rect 552 6480 15364 6502
rect 1397 6443 1455 6449
rect 1397 6409 1409 6443
rect 1443 6440 1455 6443
rect 1486 6440 1492 6452
rect 1443 6412 1492 6440
rect 1443 6409 1455 6412
rect 1397 6403 1455 6409
rect 1486 6400 1492 6412
rect 1544 6400 1550 6452
rect 1949 6443 2007 6449
rect 1949 6409 1961 6443
rect 1995 6440 2007 6443
rect 2130 6440 2136 6452
rect 1995 6412 2136 6440
rect 1995 6409 2007 6412
rect 1949 6403 2007 6409
rect 2130 6400 2136 6412
rect 2188 6400 2194 6452
rect 2409 6443 2467 6449
rect 2409 6409 2421 6443
rect 2455 6440 2467 6443
rect 2590 6440 2596 6452
rect 2455 6412 2596 6440
rect 2455 6409 2467 6412
rect 2409 6403 2467 6409
rect 2590 6400 2596 6412
rect 2648 6400 2654 6452
rect 2777 6443 2835 6449
rect 2777 6409 2789 6443
rect 2823 6440 2835 6443
rect 2958 6440 2964 6452
rect 2823 6412 2964 6440
rect 2823 6409 2835 6412
rect 2777 6403 2835 6409
rect 2958 6400 2964 6412
rect 3016 6400 3022 6452
rect 3326 6400 3332 6452
rect 3384 6400 3390 6452
rect 3881 6443 3939 6449
rect 3881 6409 3893 6443
rect 3927 6440 3939 6443
rect 4062 6440 4068 6452
rect 3927 6412 4068 6440
rect 3927 6409 3939 6412
rect 3881 6403 3939 6409
rect 4062 6400 4068 6412
rect 4120 6400 4126 6452
rect 4430 6400 4436 6452
rect 4488 6440 4494 6452
rect 4525 6443 4583 6449
rect 4525 6440 4537 6443
rect 4488 6412 4537 6440
rect 4488 6400 4494 6412
rect 4525 6409 4537 6412
rect 4571 6409 4583 6443
rect 4525 6403 4583 6409
rect 4798 6400 4804 6452
rect 4856 6400 4862 6452
rect 5169 6443 5227 6449
rect 5169 6409 5181 6443
rect 5215 6440 5227 6443
rect 5442 6440 5448 6452
rect 5215 6412 5448 6440
rect 5215 6409 5227 6412
rect 5169 6403 5227 6409
rect 5442 6400 5448 6412
rect 5500 6400 5506 6452
rect 5810 6400 5816 6452
rect 5868 6440 5874 6452
rect 5905 6443 5963 6449
rect 5905 6440 5917 6443
rect 5868 6412 5917 6440
rect 5868 6400 5874 6412
rect 5905 6409 5917 6412
rect 5951 6409 5963 6443
rect 5905 6403 5963 6409
rect 6270 6400 6276 6452
rect 6328 6440 6334 6452
rect 6365 6443 6423 6449
rect 6365 6440 6377 6443
rect 6328 6412 6377 6440
rect 6328 6400 6334 6412
rect 6365 6409 6377 6412
rect 6411 6409 6423 6443
rect 6365 6403 6423 6409
rect 6638 6400 6644 6452
rect 6696 6400 6702 6452
rect 7006 6400 7012 6452
rect 7064 6440 7070 6452
rect 7193 6443 7251 6449
rect 7193 6440 7205 6443
rect 7064 6412 7205 6440
rect 7064 6400 7070 6412
rect 7193 6409 7205 6412
rect 7239 6409 7251 6443
rect 7193 6403 7251 6409
rect 7374 6400 7380 6452
rect 7432 6440 7438 6452
rect 7653 6443 7711 6449
rect 7653 6440 7665 6443
rect 7432 6412 7665 6440
rect 7432 6400 7438 6412
rect 7653 6409 7665 6412
rect 7699 6409 7711 6443
rect 7653 6403 7711 6409
rect 7742 6400 7748 6452
rect 7800 6440 7806 6452
rect 9217 6443 9275 6449
rect 9217 6440 9229 6443
rect 7800 6412 9229 6440
rect 7800 6400 7806 6412
rect 9217 6409 9229 6412
rect 9263 6409 9275 6443
rect 9217 6403 9275 6409
rect 11974 6400 11980 6452
rect 12032 6440 12038 6452
rect 12069 6443 12127 6449
rect 12069 6440 12081 6443
rect 12032 6412 12081 6440
rect 12032 6400 12038 6412
rect 12069 6409 12081 6412
rect 12115 6409 12127 6443
rect 12069 6403 12127 6409
rect 4249 6375 4307 6381
rect 4249 6341 4261 6375
rect 4295 6341 4307 6375
rect 4816 6372 4844 6400
rect 5537 6375 5595 6381
rect 5537 6372 5549 6375
rect 4816 6344 5549 6372
rect 4249 6335 4307 6341
rect 5537 6341 5549 6344
rect 5583 6341 5595 6375
rect 5537 6335 5595 6341
rect 4264 6304 4292 6335
rect 8846 6332 8852 6384
rect 8904 6332 8910 6384
rect 8938 6332 8944 6384
rect 8996 6372 9002 6384
rect 9677 6375 9735 6381
rect 9677 6372 9689 6375
rect 8996 6344 9689 6372
rect 8996 6332 9002 6344
rect 9677 6341 9689 6344
rect 9723 6341 9735 6375
rect 9677 6335 9735 6341
rect 13817 6375 13875 6381
rect 13817 6341 13829 6375
rect 13863 6372 13875 6375
rect 14274 6372 14280 6384
rect 13863 6344 14280 6372
rect 13863 6341 13875 6344
rect 13817 6335 13875 6341
rect 14274 6332 14280 6344
rect 14332 6332 14338 6384
rect 5166 6304 5172 6316
rect 4264 6276 5172 6304
rect 5166 6264 5172 6276
rect 5224 6264 5230 6316
rect 8478 6264 8484 6316
rect 8536 6304 8542 6316
rect 8757 6307 8815 6313
rect 8757 6304 8769 6307
rect 8536 6276 8769 6304
rect 8536 6264 8542 6276
rect 8757 6273 8769 6276
rect 8803 6273 8815 6307
rect 8864 6304 8892 6332
rect 11057 6307 11115 6313
rect 11057 6304 11069 6307
rect 8864 6276 11069 6304
rect 8757 6267 8815 6273
rect 11057 6273 11069 6276
rect 11103 6273 11115 6307
rect 11057 6267 11115 6273
rect 12618 6264 12624 6316
rect 12676 6264 12682 6316
rect 13538 6264 13544 6316
rect 13596 6304 13602 6316
rect 14642 6304 14648 6316
rect 13596 6276 14648 6304
rect 13596 6264 13602 6276
rect 14642 6264 14648 6276
rect 14700 6264 14706 6316
rect 750 6196 756 6248
rect 808 6236 814 6248
rect 1121 6239 1179 6245
rect 1121 6236 1133 6239
rect 808 6208 1133 6236
rect 808 6196 814 6208
rect 1121 6205 1133 6208
rect 1167 6236 1179 6239
rect 1302 6236 1308 6248
rect 1167 6208 1308 6236
rect 1167 6205 1179 6208
rect 1121 6199 1179 6205
rect 1302 6196 1308 6208
rect 1360 6236 1366 6248
rect 1765 6239 1823 6245
rect 1765 6236 1777 6239
rect 1360 6208 1777 6236
rect 1360 6196 1366 6208
rect 1765 6205 1777 6208
rect 1811 6236 1823 6239
rect 2225 6239 2283 6245
rect 2225 6236 2237 6239
rect 1811 6208 2237 6236
rect 1811 6205 1823 6208
rect 1765 6199 1823 6205
rect 2225 6205 2237 6208
rect 2271 6236 2283 6239
rect 2593 6239 2651 6245
rect 2593 6236 2605 6239
rect 2271 6208 2605 6236
rect 2271 6205 2283 6208
rect 2225 6199 2283 6205
rect 2593 6205 2605 6208
rect 2639 6236 2651 6239
rect 3513 6239 3571 6245
rect 3513 6236 3525 6239
rect 2639 6208 3525 6236
rect 2639 6205 2651 6208
rect 2593 6199 2651 6205
rect 3513 6205 3525 6208
rect 3559 6205 3571 6239
rect 3513 6199 3571 6205
rect 3528 6168 3556 6199
rect 3602 6196 3608 6248
rect 3660 6236 3666 6248
rect 3697 6239 3755 6245
rect 3697 6236 3709 6239
rect 3660 6208 3709 6236
rect 3660 6196 3666 6208
rect 3697 6205 3709 6208
rect 3743 6205 3755 6239
rect 3697 6199 3755 6205
rect 3878 6196 3884 6248
rect 3936 6236 3942 6248
rect 4065 6239 4123 6245
rect 4065 6236 4077 6239
rect 3936 6208 4077 6236
rect 3936 6196 3942 6208
rect 4065 6205 4077 6208
rect 4111 6205 4123 6239
rect 4065 6199 4123 6205
rect 4522 6196 4528 6248
rect 4580 6196 4586 6248
rect 4706 6196 4712 6248
rect 4764 6196 4770 6248
rect 5350 6196 5356 6248
rect 5408 6196 5414 6248
rect 6089 6239 6147 6245
rect 6089 6205 6101 6239
rect 6135 6205 6147 6239
rect 6089 6199 6147 6205
rect 4540 6168 4568 6196
rect 3528 6140 4568 6168
rect 4893 6171 4951 6177
rect 4893 6137 4905 6171
rect 4939 6168 4951 6171
rect 4982 6168 4988 6180
rect 4939 6140 4988 6168
rect 4939 6137 4951 6140
rect 4893 6131 4951 6137
rect 4982 6128 4988 6140
rect 5040 6128 5046 6180
rect 6104 6168 6132 6199
rect 6178 6196 6184 6248
rect 6236 6196 6242 6248
rect 6822 6196 6828 6248
rect 6880 6196 6886 6248
rect 7374 6196 7380 6248
rect 7432 6196 7438 6248
rect 7837 6239 7895 6245
rect 7837 6205 7849 6239
rect 7883 6236 7895 6239
rect 8846 6236 8852 6248
rect 7883 6208 8852 6236
rect 7883 6205 7895 6208
rect 7837 6199 7895 6205
rect 8846 6196 8852 6208
rect 8904 6196 8910 6248
rect 9033 6239 9091 6245
rect 9033 6205 9045 6239
rect 9079 6205 9091 6239
rect 9033 6199 9091 6205
rect 6914 6168 6920 6180
rect 6104 6140 6920 6168
rect 6914 6128 6920 6140
rect 6972 6128 6978 6180
rect 9048 6100 9076 6199
rect 9398 6196 9404 6248
rect 9456 6236 9462 6248
rect 9861 6239 9919 6245
rect 9861 6236 9873 6239
rect 9456 6208 9873 6236
rect 9456 6196 9462 6208
rect 9861 6205 9873 6208
rect 9907 6205 9919 6239
rect 9861 6199 9919 6205
rect 10042 6196 10048 6248
rect 10100 6236 10106 6248
rect 10229 6239 10287 6245
rect 10229 6236 10241 6239
rect 10100 6208 10241 6236
rect 10100 6196 10106 6208
rect 10229 6205 10241 6208
rect 10275 6205 10287 6239
rect 10229 6199 10287 6205
rect 10318 6196 10324 6248
rect 10376 6236 10382 6248
rect 10597 6239 10655 6245
rect 10597 6236 10609 6239
rect 10376 6208 10609 6236
rect 10376 6196 10382 6208
rect 10597 6205 10609 6208
rect 10643 6205 10655 6239
rect 10597 6199 10655 6205
rect 11609 6239 11667 6245
rect 11609 6205 11621 6239
rect 11655 6236 11667 6239
rect 11882 6236 11888 6248
rect 11655 6208 11888 6236
rect 11655 6205 11667 6208
rect 11609 6199 11667 6205
rect 11882 6196 11888 6208
rect 11940 6196 11946 6248
rect 13998 6196 14004 6248
rect 14056 6196 14062 6248
rect 9493 6171 9551 6177
rect 9493 6137 9505 6171
rect 9539 6168 9551 6171
rect 10962 6168 10968 6180
rect 9539 6140 10968 6168
rect 9539 6137 9551 6140
rect 9493 6131 9551 6137
rect 10962 6128 10968 6140
rect 11020 6128 11026 6180
rect 12342 6128 12348 6180
rect 12400 6128 12406 6180
rect 14182 6128 14188 6180
rect 14240 6168 14246 6180
rect 14553 6171 14611 6177
rect 14553 6168 14565 6171
rect 14240 6140 14565 6168
rect 14240 6128 14246 6140
rect 14553 6137 14565 6140
rect 14599 6137 14611 6171
rect 14553 6131 14611 6137
rect 9950 6100 9956 6112
rect 9048 6072 9956 6100
rect 9950 6060 9956 6072
rect 10008 6060 10014 6112
rect 10042 6060 10048 6112
rect 10100 6060 10106 6112
rect 10410 6060 10416 6112
rect 10468 6060 10474 6112
rect 12802 6060 12808 6112
rect 12860 6060 12866 6112
rect 12897 6103 12955 6109
rect 12897 6069 12909 6103
rect 12943 6100 12955 6103
rect 12986 6100 12992 6112
rect 12943 6072 12992 6100
rect 12943 6069 12955 6072
rect 12897 6063 12955 6069
rect 12986 6060 12992 6072
rect 13044 6060 13050 6112
rect 13265 6103 13323 6109
rect 13265 6069 13277 6103
rect 13311 6100 13323 6103
rect 13814 6100 13820 6112
rect 13311 6072 13820 6100
rect 13311 6069 13323 6072
rect 13265 6063 13323 6069
rect 13814 6060 13820 6072
rect 13872 6060 13878 6112
rect 14090 6060 14096 6112
rect 14148 6060 14154 6112
rect 14461 6103 14519 6109
rect 14461 6069 14473 6103
rect 14507 6100 14519 6103
rect 14826 6100 14832 6112
rect 14507 6072 14832 6100
rect 14507 6069 14519 6072
rect 14461 6063 14519 6069
rect 14826 6060 14832 6072
rect 14884 6060 14890 6112
rect 552 6010 15520 6032
rect 552 5958 4100 6010
rect 4152 5958 4164 6010
rect 4216 5958 4228 6010
rect 4280 5958 4292 6010
rect 4344 5958 4356 6010
rect 4408 5958 7802 6010
rect 7854 5958 7866 6010
rect 7918 5958 7930 6010
rect 7982 5958 7994 6010
rect 8046 5958 8058 6010
rect 8110 5958 11504 6010
rect 11556 5958 11568 6010
rect 11620 5958 11632 6010
rect 11684 5958 11696 6010
rect 11748 5958 11760 6010
rect 11812 5958 15206 6010
rect 15258 5958 15270 6010
rect 15322 5958 15334 6010
rect 15386 5958 15398 6010
rect 15450 5958 15462 6010
rect 15514 5958 15520 6010
rect 552 5936 15520 5958
rect 1118 5856 1124 5908
rect 1176 5856 1182 5908
rect 1581 5899 1639 5905
rect 1581 5865 1593 5899
rect 1627 5896 1639 5899
rect 1854 5896 1860 5908
rect 1627 5868 1860 5896
rect 1627 5865 1639 5868
rect 1581 5859 1639 5865
rect 1854 5856 1860 5868
rect 1912 5856 1918 5908
rect 3694 5856 3700 5908
rect 3752 5896 3758 5908
rect 3973 5899 4031 5905
rect 3973 5896 3985 5899
rect 3752 5868 3985 5896
rect 3752 5856 3758 5868
rect 3973 5865 3985 5868
rect 4019 5865 4031 5899
rect 3973 5859 4031 5865
rect 5626 5856 5632 5908
rect 5684 5856 5690 5908
rect 6733 5899 6791 5905
rect 6733 5865 6745 5899
rect 6779 5896 6791 5899
rect 6822 5896 6828 5908
rect 6779 5868 6828 5896
rect 6779 5865 6791 5868
rect 6733 5859 6791 5865
rect 6822 5856 6828 5868
rect 6880 5856 6886 5908
rect 7098 5856 7104 5908
rect 7156 5856 7162 5908
rect 7190 5856 7196 5908
rect 7248 5896 7254 5908
rect 8938 5896 8944 5908
rect 7248 5868 8944 5896
rect 7248 5856 7254 5868
rect 8938 5856 8944 5868
rect 8996 5856 9002 5908
rect 9033 5899 9091 5905
rect 9033 5865 9045 5899
rect 9079 5896 9091 5899
rect 10042 5896 10048 5908
rect 9079 5868 10048 5896
rect 9079 5865 9091 5868
rect 9033 5859 9091 5865
rect 10042 5856 10048 5868
rect 10100 5856 10106 5908
rect 10686 5856 10692 5908
rect 10744 5856 10750 5908
rect 10962 5856 10968 5908
rect 11020 5856 11026 5908
rect 11793 5899 11851 5905
rect 11793 5865 11805 5899
rect 11839 5896 11851 5899
rect 11882 5896 11888 5908
rect 11839 5868 11888 5896
rect 11839 5865 11851 5868
rect 11793 5859 11851 5865
rect 11882 5856 11888 5868
rect 11940 5856 11946 5908
rect 12161 5899 12219 5905
rect 12161 5865 12173 5899
rect 12207 5896 12219 5899
rect 12250 5896 12256 5908
rect 12207 5868 12256 5896
rect 12207 5865 12219 5868
rect 12161 5859 12219 5865
rect 12250 5856 12256 5868
rect 12308 5896 12314 5908
rect 14826 5896 14832 5908
rect 12308 5868 14832 5896
rect 12308 5856 12314 5868
rect 14826 5856 14832 5868
rect 14884 5856 14890 5908
rect 3234 5788 3240 5840
rect 3292 5788 3298 5840
rect 6273 5831 6331 5837
rect 4540 5800 6040 5828
rect 1302 5720 1308 5772
rect 1360 5760 1366 5772
rect 1397 5763 1455 5769
rect 1397 5760 1409 5763
rect 1360 5732 1409 5760
rect 1360 5720 1366 5732
rect 1397 5729 1409 5732
rect 1443 5729 1455 5763
rect 1397 5723 1455 5729
rect 3510 5720 3516 5772
rect 3568 5720 3574 5772
rect 3789 5695 3847 5701
rect 3789 5661 3801 5695
rect 3835 5692 3847 5695
rect 4540 5692 4568 5800
rect 4614 5720 4620 5772
rect 4672 5760 4678 5772
rect 5261 5763 5319 5769
rect 5261 5760 5273 5763
rect 4672 5732 5273 5760
rect 4672 5720 4678 5732
rect 5261 5729 5273 5732
rect 5307 5729 5319 5763
rect 5261 5723 5319 5729
rect 4890 5692 4896 5704
rect 3835 5664 4896 5692
rect 3835 5661 3847 5664
rect 3789 5655 3847 5661
rect 4890 5652 4896 5664
rect 4948 5652 4954 5704
rect 5077 5695 5135 5701
rect 5077 5661 5089 5695
rect 5123 5661 5135 5695
rect 5077 5655 5135 5661
rect 5169 5695 5227 5701
rect 5169 5661 5181 5695
rect 5215 5661 5227 5695
rect 6012 5692 6040 5800
rect 6273 5797 6285 5831
rect 6319 5828 6331 5831
rect 10137 5831 10195 5837
rect 6319 5800 8248 5828
rect 6319 5797 6331 5800
rect 6273 5791 6331 5797
rect 6365 5763 6423 5769
rect 6365 5729 6377 5763
rect 6411 5760 6423 5763
rect 7193 5763 7251 5769
rect 7193 5760 7205 5763
rect 6411 5732 7205 5760
rect 6411 5729 6423 5732
rect 6365 5723 6423 5729
rect 7193 5729 7205 5732
rect 7239 5760 7251 5763
rect 7650 5760 7656 5772
rect 7239 5732 7656 5760
rect 7239 5729 7251 5732
rect 7193 5723 7251 5729
rect 7650 5720 7656 5732
rect 7708 5720 7714 5772
rect 8220 5769 8248 5800
rect 10137 5797 10149 5831
rect 10183 5828 10195 5831
rect 10318 5828 10324 5840
rect 10183 5800 10324 5828
rect 10183 5797 10195 5800
rect 10137 5791 10195 5797
rect 10318 5788 10324 5800
rect 10376 5788 10382 5840
rect 8205 5763 8263 5769
rect 8205 5729 8217 5763
rect 8251 5760 8263 5763
rect 8570 5760 8576 5772
rect 8251 5732 8576 5760
rect 8251 5729 8263 5732
rect 8205 5723 8263 5729
rect 8570 5720 8576 5732
rect 8628 5720 8634 5772
rect 8846 5720 8852 5772
rect 8904 5720 8910 5772
rect 8941 5763 8999 5769
rect 8941 5729 8953 5763
rect 8987 5760 8999 5763
rect 9306 5760 9312 5772
rect 8987 5732 9312 5760
rect 8987 5729 8999 5732
rect 8941 5723 8999 5729
rect 9306 5720 9312 5732
rect 9364 5720 9370 5772
rect 10704 5760 10732 5856
rect 10870 5788 10876 5840
rect 10928 5828 10934 5840
rect 12805 5831 12863 5837
rect 12805 5828 12817 5831
rect 10928 5800 12817 5828
rect 10928 5788 10934 5800
rect 12805 5797 12817 5800
rect 12851 5797 12863 5831
rect 12805 5791 12863 5797
rect 13814 5788 13820 5840
rect 13872 5828 13878 5840
rect 13872 5800 14412 5828
rect 13872 5788 13878 5800
rect 10781 5763 10839 5769
rect 10781 5760 10793 5763
rect 10152 5732 10364 5760
rect 10704 5732 10793 5760
rect 6089 5695 6147 5701
rect 6089 5692 6101 5695
rect 6012 5664 6101 5692
rect 5169 5655 5227 5661
rect 6089 5661 6101 5664
rect 6135 5661 6147 5695
rect 6089 5655 6147 5661
rect 2869 5627 2927 5633
rect 2869 5593 2881 5627
rect 2915 5624 2927 5627
rect 3050 5624 3056 5636
rect 2915 5596 3056 5624
rect 2915 5593 2927 5596
rect 2869 5587 2927 5593
rect 3050 5584 3056 5596
rect 3108 5584 3114 5636
rect 3421 5627 3479 5633
rect 3421 5593 3433 5627
rect 3467 5624 3479 5627
rect 3605 5627 3663 5633
rect 3605 5624 3617 5627
rect 3467 5596 3617 5624
rect 3467 5593 3479 5596
rect 3421 5587 3479 5593
rect 3605 5593 3617 5596
rect 3651 5593 3663 5627
rect 3605 5587 3663 5593
rect 2958 5516 2964 5568
rect 3016 5556 3022 5568
rect 3237 5559 3295 5565
rect 3237 5556 3249 5559
rect 3016 5528 3249 5556
rect 3016 5516 3022 5528
rect 3237 5525 3249 5528
rect 3283 5525 3295 5559
rect 5092 5556 5120 5655
rect 5184 5624 5212 5655
rect 6730 5652 6736 5704
rect 6788 5692 6794 5704
rect 7009 5695 7067 5701
rect 7009 5692 7021 5695
rect 6788 5664 7021 5692
rect 6788 5652 6794 5664
rect 7009 5661 7021 5664
rect 7055 5692 7067 5695
rect 7466 5692 7472 5704
rect 7055 5664 7472 5692
rect 7055 5661 7067 5664
rect 7009 5655 7067 5661
rect 7466 5652 7472 5664
rect 7524 5652 7530 5704
rect 8481 5695 8539 5701
rect 8481 5661 8493 5695
rect 8527 5692 8539 5695
rect 8527 5664 8616 5692
rect 8527 5661 8539 5664
rect 8481 5655 8539 5661
rect 8588 5633 8616 5664
rect 8573 5627 8631 5633
rect 5184 5596 7696 5624
rect 6730 5556 6736 5568
rect 5092 5528 6736 5556
rect 3237 5519 3295 5525
rect 6730 5516 6736 5528
rect 6788 5516 6794 5568
rect 7558 5516 7564 5568
rect 7616 5516 7622 5568
rect 7668 5556 7696 5596
rect 8573 5593 8585 5627
rect 8619 5593 8631 5627
rect 8864 5624 8892 5720
rect 9217 5695 9275 5701
rect 9217 5661 9229 5695
rect 9263 5692 9275 5695
rect 9398 5692 9404 5704
rect 9263 5664 9404 5692
rect 9263 5661 9275 5664
rect 9217 5655 9275 5661
rect 9398 5652 9404 5664
rect 9456 5652 9462 5704
rect 9490 5652 9496 5704
rect 9548 5692 9554 5704
rect 10152 5692 10180 5732
rect 9548 5664 10180 5692
rect 9548 5652 9554 5664
rect 10226 5652 10232 5704
rect 10284 5652 10290 5704
rect 10336 5701 10364 5732
rect 10781 5729 10793 5732
rect 10827 5729 10839 5763
rect 10781 5723 10839 5729
rect 11330 5720 11336 5772
rect 11388 5720 11394 5772
rect 11425 5763 11483 5769
rect 11425 5729 11437 5763
rect 11471 5760 11483 5763
rect 11471 5732 12572 5760
rect 11471 5729 11483 5732
rect 11425 5723 11483 5729
rect 12544 5704 12572 5732
rect 12710 5720 12716 5772
rect 12768 5760 12774 5772
rect 13357 5763 13415 5769
rect 13357 5760 13369 5763
rect 12768 5732 13369 5760
rect 12768 5720 12774 5732
rect 13357 5729 13369 5732
rect 13403 5760 13415 5763
rect 13538 5760 13544 5772
rect 13403 5732 13544 5760
rect 13403 5729 13415 5732
rect 13357 5723 13415 5729
rect 13538 5720 13544 5732
rect 13596 5720 13602 5772
rect 13906 5720 13912 5772
rect 13964 5720 13970 5772
rect 14384 5769 14412 5800
rect 14369 5763 14427 5769
rect 14369 5729 14381 5763
rect 14415 5729 14427 5763
rect 14369 5723 14427 5729
rect 10321 5695 10379 5701
rect 10321 5661 10333 5695
rect 10367 5692 10379 5695
rect 11146 5692 11152 5704
rect 10367 5664 11152 5692
rect 10367 5661 10379 5664
rect 10321 5655 10379 5661
rect 11146 5652 11152 5664
rect 11204 5652 11210 5704
rect 11517 5695 11575 5701
rect 11517 5661 11529 5695
rect 11563 5661 11575 5695
rect 11517 5655 11575 5661
rect 9769 5627 9827 5633
rect 9769 5624 9781 5627
rect 8864 5596 9781 5624
rect 8573 5587 8631 5593
rect 9769 5593 9781 5596
rect 9815 5593 9827 5627
rect 9769 5587 9827 5593
rect 10134 5584 10140 5636
rect 10192 5624 10198 5636
rect 11532 5624 11560 5655
rect 11974 5652 11980 5704
rect 12032 5692 12038 5704
rect 12253 5695 12311 5701
rect 12253 5692 12265 5695
rect 12032 5664 12265 5692
rect 12032 5652 12038 5664
rect 12253 5661 12265 5664
rect 12299 5661 12311 5695
rect 12253 5655 12311 5661
rect 12345 5695 12403 5701
rect 12345 5661 12357 5695
rect 12391 5661 12403 5695
rect 12345 5655 12403 5661
rect 12360 5624 12388 5655
rect 12526 5652 12532 5704
rect 12584 5652 12590 5704
rect 13998 5652 14004 5704
rect 14056 5652 14062 5704
rect 14093 5695 14151 5701
rect 14093 5661 14105 5695
rect 14139 5661 14151 5695
rect 14093 5655 14151 5661
rect 12618 5624 12624 5636
rect 10192 5596 12624 5624
rect 10192 5584 10198 5596
rect 12618 5584 12624 5596
rect 12676 5584 12682 5636
rect 12894 5584 12900 5636
rect 12952 5624 12958 5636
rect 14108 5624 14136 5655
rect 14550 5652 14556 5704
rect 14608 5652 14614 5704
rect 12952 5596 14136 5624
rect 12952 5584 12958 5596
rect 10597 5559 10655 5565
rect 10597 5556 10609 5559
rect 7668 5528 10609 5556
rect 10597 5525 10609 5528
rect 10643 5525 10655 5559
rect 10597 5519 10655 5525
rect 11238 5516 11244 5568
rect 11296 5556 11302 5568
rect 12250 5556 12256 5568
rect 11296 5528 12256 5556
rect 11296 5516 11302 5528
rect 12250 5516 12256 5528
rect 12308 5516 12314 5568
rect 13541 5559 13599 5565
rect 13541 5525 13553 5559
rect 13587 5556 13599 5559
rect 13722 5556 13728 5568
rect 13587 5528 13728 5556
rect 13587 5525 13599 5528
rect 13541 5519 13599 5525
rect 13722 5516 13728 5528
rect 13780 5516 13786 5568
rect 552 5466 15364 5488
rect 552 5414 2249 5466
rect 2301 5414 2313 5466
rect 2365 5414 2377 5466
rect 2429 5414 2441 5466
rect 2493 5414 2505 5466
rect 2557 5414 5951 5466
rect 6003 5414 6015 5466
rect 6067 5414 6079 5466
rect 6131 5414 6143 5466
rect 6195 5414 6207 5466
rect 6259 5414 9653 5466
rect 9705 5414 9717 5466
rect 9769 5414 9781 5466
rect 9833 5414 9845 5466
rect 9897 5414 9909 5466
rect 9961 5414 13355 5466
rect 13407 5414 13419 5466
rect 13471 5414 13483 5466
rect 13535 5414 13547 5466
rect 13599 5414 13611 5466
rect 13663 5414 15364 5466
rect 552 5392 15364 5414
rect 4706 5312 4712 5364
rect 4764 5352 4770 5364
rect 4801 5355 4859 5361
rect 4801 5352 4813 5355
rect 4764 5324 4813 5352
rect 4764 5312 4770 5324
rect 4801 5321 4813 5324
rect 4847 5321 4859 5355
rect 4801 5315 4859 5321
rect 5166 5312 5172 5364
rect 5224 5352 5230 5364
rect 9306 5352 9312 5364
rect 5224 5324 9312 5352
rect 5224 5312 5230 5324
rect 9306 5312 9312 5324
rect 9364 5312 9370 5364
rect 10594 5312 10600 5364
rect 10652 5352 10658 5364
rect 10965 5355 11023 5361
rect 10965 5352 10977 5355
rect 10652 5324 10977 5352
rect 10652 5312 10658 5324
rect 10965 5321 10977 5324
rect 11011 5321 11023 5355
rect 10965 5315 11023 5321
rect 11146 5312 11152 5364
rect 11204 5352 11210 5364
rect 11333 5355 11391 5361
rect 11333 5352 11345 5355
rect 11204 5324 11345 5352
rect 11204 5312 11210 5324
rect 11333 5321 11345 5324
rect 11379 5321 11391 5355
rect 11333 5315 11391 5321
rect 11514 5312 11520 5364
rect 11572 5352 11578 5364
rect 12253 5355 12311 5361
rect 11572 5324 11836 5352
rect 11572 5312 11578 5324
rect 8846 5244 8852 5296
rect 8904 5284 8910 5296
rect 11609 5287 11667 5293
rect 11609 5284 11621 5287
rect 8904 5256 11621 5284
rect 8904 5244 8910 5256
rect 11609 5253 11621 5256
rect 11655 5253 11667 5287
rect 11609 5247 11667 5253
rect 5442 5176 5448 5228
rect 5500 5176 5506 5228
rect 5626 5176 5632 5228
rect 5684 5216 5690 5228
rect 8938 5216 8944 5228
rect 5684 5188 6040 5216
rect 5684 5176 5690 5188
rect 2317 5151 2375 5157
rect 2317 5117 2329 5151
rect 2363 5117 2375 5151
rect 2317 5111 2375 5117
rect 2593 5151 2651 5157
rect 2593 5117 2605 5151
rect 2639 5117 2651 5151
rect 2593 5111 2651 5117
rect 2777 5151 2835 5157
rect 2777 5117 2789 5151
rect 2823 5148 2835 5151
rect 2961 5151 3019 5157
rect 2961 5148 2973 5151
rect 2823 5120 2973 5148
rect 2823 5117 2835 5120
rect 2777 5111 2835 5117
rect 2961 5117 2973 5120
rect 3007 5117 3019 5151
rect 2961 5111 3019 5117
rect 2130 4972 2136 5024
rect 2188 4972 2194 5024
rect 2332 5012 2360 5111
rect 2608 5080 2636 5111
rect 3050 5108 3056 5160
rect 3108 5148 3114 5160
rect 3694 5148 3700 5160
rect 3108 5120 3700 5148
rect 3108 5108 3114 5120
rect 3694 5108 3700 5120
rect 3752 5108 3758 5160
rect 4706 5108 4712 5160
rect 4764 5148 4770 5160
rect 5166 5148 5172 5160
rect 4764 5120 5172 5148
rect 4764 5108 4770 5120
rect 5166 5108 5172 5120
rect 5224 5108 5230 5160
rect 6012 5157 6040 5188
rect 6748 5188 8944 5216
rect 6748 5157 6776 5188
rect 8938 5176 8944 5188
rect 8996 5216 9002 5228
rect 9490 5216 9496 5228
rect 8996 5188 9496 5216
rect 8996 5176 9002 5188
rect 9490 5176 9496 5188
rect 9548 5176 9554 5228
rect 10137 5219 10195 5225
rect 10137 5216 10149 5219
rect 9646 5188 10149 5216
rect 5997 5151 6055 5157
rect 5997 5117 6009 5151
rect 6043 5117 6055 5151
rect 5997 5111 6055 5117
rect 6733 5151 6791 5157
rect 6733 5117 6745 5151
rect 6779 5117 6791 5151
rect 6733 5111 6791 5117
rect 7377 5151 7435 5157
rect 7377 5117 7389 5151
rect 7423 5148 7435 5151
rect 7558 5148 7564 5160
rect 7423 5120 7564 5148
rect 7423 5117 7435 5120
rect 7377 5111 7435 5117
rect 7558 5108 7564 5120
rect 7616 5108 7622 5160
rect 8570 5108 8576 5160
rect 8628 5148 8634 5160
rect 9122 5148 9128 5160
rect 8628 5120 9128 5148
rect 8628 5108 8634 5120
rect 9122 5108 9128 5120
rect 9180 5108 9186 5160
rect 9398 5108 9404 5160
rect 9456 5148 9462 5160
rect 9646 5148 9674 5188
rect 10137 5185 10149 5188
rect 10183 5216 10195 5219
rect 10183 5188 11008 5216
rect 10183 5185 10195 5188
rect 10137 5179 10195 5185
rect 10781 5151 10839 5157
rect 10781 5148 10793 5151
rect 9456 5120 9674 5148
rect 10704 5120 10793 5148
rect 9456 5108 9462 5120
rect 2682 5080 2688 5092
rect 2608 5052 2688 5080
rect 2682 5040 2688 5052
rect 2740 5080 2746 5092
rect 4246 5080 4252 5092
rect 2740 5052 4252 5080
rect 2740 5040 2746 5052
rect 4246 5040 4252 5052
rect 4304 5040 4310 5092
rect 4430 5040 4436 5092
rect 4488 5080 4494 5092
rect 7193 5083 7251 5089
rect 7193 5080 7205 5083
rect 4488 5052 7205 5080
rect 4488 5040 4494 5052
rect 7193 5049 7205 5052
rect 7239 5080 7251 5083
rect 7282 5080 7288 5092
rect 7239 5052 7288 5080
rect 7239 5049 7251 5052
rect 7193 5043 7251 5049
rect 7282 5040 7288 5052
rect 7340 5040 7346 5092
rect 8202 5040 8208 5092
rect 8260 5080 8266 5092
rect 10134 5080 10140 5092
rect 8260 5052 10140 5080
rect 8260 5040 8266 5052
rect 10134 5040 10140 5052
rect 10192 5040 10198 5092
rect 10226 5040 10232 5092
rect 10284 5080 10290 5092
rect 10284 5052 10548 5080
rect 10284 5040 10290 5052
rect 10520 5024 10548 5052
rect 2958 5012 2964 5024
rect 2332 4984 2964 5012
rect 2958 4972 2964 4984
rect 3016 4972 3022 5024
rect 5258 4972 5264 5024
rect 5316 4972 5322 5024
rect 5534 4972 5540 5024
rect 5592 5012 5598 5024
rect 5813 5015 5871 5021
rect 5813 5012 5825 5015
rect 5592 4984 5825 5012
rect 5592 4972 5598 4984
rect 5813 4981 5825 4984
rect 5859 4981 5871 5015
rect 5813 4975 5871 4981
rect 6178 4972 6184 5024
rect 6236 5012 6242 5024
rect 6641 5015 6699 5021
rect 6641 5012 6653 5015
rect 6236 4984 6653 5012
rect 6236 4972 6242 4984
rect 6641 4981 6653 4984
rect 6687 5012 6699 5015
rect 9490 5012 9496 5024
rect 6687 4984 9496 5012
rect 6687 4981 6699 4984
rect 6641 4975 6699 4981
rect 9490 4972 9496 4984
rect 9548 4972 9554 5024
rect 10318 4972 10324 5024
rect 10376 4972 10382 5024
rect 10502 4972 10508 5024
rect 10560 4972 10566 5024
rect 10704 5021 10732 5120
rect 10781 5117 10793 5120
rect 10827 5117 10839 5151
rect 10781 5111 10839 5117
rect 10980 5080 11008 5188
rect 11054 5176 11060 5228
rect 11112 5216 11118 5228
rect 11808 5216 11836 5324
rect 12253 5321 12265 5355
rect 12299 5352 12311 5355
rect 12342 5352 12348 5364
rect 12299 5324 12348 5352
rect 12299 5321 12311 5324
rect 12253 5315 12311 5321
rect 12342 5312 12348 5324
rect 12400 5312 12406 5364
rect 12526 5312 12532 5364
rect 12584 5352 12590 5364
rect 12584 5324 14320 5352
rect 12584 5312 12590 5324
rect 12618 5216 12624 5228
rect 11112 5188 11652 5216
rect 11808 5188 12112 5216
rect 11112 5176 11118 5188
rect 11422 5108 11428 5160
rect 11480 5148 11486 5160
rect 11517 5151 11575 5157
rect 11517 5148 11529 5151
rect 11480 5120 11529 5148
rect 11480 5108 11486 5120
rect 11517 5117 11529 5120
rect 11563 5117 11575 5151
rect 11624 5148 11652 5188
rect 12084 5157 12112 5188
rect 12176 5188 12624 5216
rect 12176 5160 12204 5188
rect 12618 5176 12624 5188
rect 12676 5216 12682 5228
rect 12805 5219 12863 5225
rect 12805 5216 12817 5219
rect 12676 5188 12817 5216
rect 12676 5176 12682 5188
rect 12805 5185 12817 5188
rect 12851 5185 12863 5219
rect 12805 5179 12863 5185
rect 14001 5219 14059 5225
rect 14001 5185 14013 5219
rect 14047 5216 14059 5219
rect 14090 5216 14096 5228
rect 14047 5188 14096 5216
rect 14047 5185 14059 5188
rect 14001 5179 14059 5185
rect 14090 5176 14096 5188
rect 14148 5176 14154 5228
rect 14292 5225 14320 5324
rect 14277 5219 14335 5225
rect 14277 5185 14289 5219
rect 14323 5216 14335 5219
rect 14918 5216 14924 5228
rect 14323 5188 14924 5216
rect 14323 5185 14335 5188
rect 14277 5179 14335 5185
rect 14918 5176 14924 5188
rect 14976 5176 14982 5228
rect 11793 5151 11851 5157
rect 11793 5148 11805 5151
rect 11624 5120 11805 5148
rect 11517 5111 11575 5117
rect 11793 5117 11805 5120
rect 11839 5117 11851 5151
rect 11793 5111 11851 5117
rect 12069 5151 12127 5157
rect 12069 5117 12081 5151
rect 12115 5117 12127 5151
rect 12069 5111 12127 5117
rect 12158 5108 12164 5160
rect 12216 5108 12222 5160
rect 12250 5108 12256 5160
rect 12308 5148 12314 5160
rect 13265 5151 13323 5157
rect 13265 5148 13277 5151
rect 12308 5120 13277 5148
rect 12308 5108 12314 5120
rect 13265 5117 13277 5120
rect 13311 5117 13323 5151
rect 13265 5111 13323 5117
rect 13633 5151 13691 5157
rect 13633 5117 13645 5151
rect 13679 5148 13691 5151
rect 13722 5148 13728 5160
rect 13679 5120 13728 5148
rect 13679 5117 13691 5120
rect 13633 5111 13691 5117
rect 13722 5108 13728 5120
rect 13780 5108 13786 5160
rect 13906 5108 13912 5160
rect 13964 5108 13970 5160
rect 12621 5083 12679 5089
rect 10980 5052 12296 5080
rect 12268 5024 12296 5052
rect 12621 5049 12633 5083
rect 12667 5080 12679 5083
rect 13924 5080 13952 5108
rect 12667 5052 13952 5080
rect 12667 5049 12679 5052
rect 12621 5043 12679 5049
rect 10689 5015 10747 5021
rect 10689 4981 10701 5015
rect 10735 4981 10747 5015
rect 10689 4975 10747 4981
rect 11054 4972 11060 5024
rect 11112 5012 11118 5024
rect 11885 5015 11943 5021
rect 11885 5012 11897 5015
rect 11112 4984 11897 5012
rect 11112 4972 11118 4984
rect 11885 4981 11897 4984
rect 11931 4981 11943 5015
rect 11885 4975 11943 4981
rect 12250 4972 12256 5024
rect 12308 4972 12314 5024
rect 12342 4972 12348 5024
rect 12400 5012 12406 5024
rect 12636 5012 12664 5043
rect 12400 4984 12664 5012
rect 12400 4972 12406 4984
rect 12710 4972 12716 5024
rect 12768 4972 12774 5024
rect 13078 4972 13084 5024
rect 13136 4972 13142 5024
rect 13725 5015 13783 5021
rect 13725 4981 13737 5015
rect 13771 5012 13783 5015
rect 13906 5012 13912 5024
rect 13771 4984 13912 5012
rect 13771 4981 13783 4984
rect 13725 4975 13783 4981
rect 13906 4972 13912 4984
rect 13964 4972 13970 5024
rect 552 4922 15520 4944
rect 552 4870 4100 4922
rect 4152 4870 4164 4922
rect 4216 4870 4228 4922
rect 4280 4870 4292 4922
rect 4344 4870 4356 4922
rect 4408 4870 7802 4922
rect 7854 4870 7866 4922
rect 7918 4870 7930 4922
rect 7982 4870 7994 4922
rect 8046 4870 8058 4922
rect 8110 4870 11504 4922
rect 11556 4870 11568 4922
rect 11620 4870 11632 4922
rect 11684 4870 11696 4922
rect 11748 4870 11760 4922
rect 11812 4870 15206 4922
rect 15258 4870 15270 4922
rect 15322 4870 15334 4922
rect 15386 4870 15398 4922
rect 15450 4870 15462 4922
rect 15514 4870 15520 4922
rect 552 4848 15520 4870
rect 2130 4768 2136 4820
rect 2188 4768 2194 4820
rect 3878 4768 3884 4820
rect 3936 4768 3942 4820
rect 4249 4811 4307 4817
rect 4249 4777 4261 4811
rect 4295 4808 4307 4811
rect 4614 4808 4620 4820
rect 4295 4780 4620 4808
rect 4295 4777 4307 4780
rect 4249 4771 4307 4777
rect 4614 4768 4620 4780
rect 4672 4768 4678 4820
rect 4890 4768 4896 4820
rect 4948 4768 4954 4820
rect 7374 4768 7380 4820
rect 7432 4768 7438 4820
rect 7837 4811 7895 4817
rect 7837 4777 7849 4811
rect 7883 4808 7895 4811
rect 9030 4808 9036 4820
rect 7883 4780 9036 4808
rect 7883 4777 7895 4780
rect 7837 4771 7895 4777
rect 9030 4768 9036 4780
rect 9088 4768 9094 4820
rect 10042 4768 10048 4820
rect 10100 4808 10106 4820
rect 10965 4811 11023 4817
rect 10965 4808 10977 4811
rect 10100 4780 10977 4808
rect 10100 4768 10106 4780
rect 10965 4777 10977 4780
rect 11011 4777 11023 4811
rect 11238 4808 11244 4820
rect 10965 4771 11023 4777
rect 11164 4780 11244 4808
rect 2148 4672 2176 4768
rect 5258 4700 5264 4752
rect 5316 4740 5322 4752
rect 8205 4743 8263 4749
rect 8205 4740 8217 4743
rect 5316 4712 8217 4740
rect 5316 4700 5322 4712
rect 8205 4709 8217 4712
rect 8251 4709 8263 4743
rect 10594 4740 10600 4752
rect 8205 4703 8263 4709
rect 10244 4712 10600 4740
rect 2317 4675 2375 4681
rect 2317 4672 2329 4675
rect 2148 4644 2329 4672
rect 2317 4641 2329 4644
rect 2363 4641 2375 4675
rect 2317 4635 2375 4641
rect 4801 4675 4859 4681
rect 4801 4641 4813 4675
rect 4847 4641 4859 4675
rect 4801 4635 4859 4641
rect 5997 4675 6055 4681
rect 5997 4641 6009 4675
rect 6043 4641 6055 4675
rect 5997 4635 6055 4641
rect 2498 4564 2504 4616
rect 2556 4564 2562 4616
rect 2593 4607 2651 4613
rect 2593 4573 2605 4607
rect 2639 4604 2651 4607
rect 3694 4604 3700 4616
rect 2639 4576 3700 4604
rect 2639 4573 2651 4576
rect 2593 4567 2651 4573
rect 3694 4564 3700 4576
rect 3752 4564 3758 4616
rect 4338 4564 4344 4616
rect 4396 4564 4402 4616
rect 4430 4564 4436 4616
rect 4488 4604 4494 4616
rect 4816 4604 4844 4635
rect 5442 4604 5448 4616
rect 4488 4576 5448 4604
rect 4488 4564 4494 4576
rect 5442 4564 5448 4576
rect 5500 4604 5506 4616
rect 5813 4607 5871 4613
rect 5813 4604 5825 4607
rect 5500 4576 5825 4604
rect 5500 4564 5506 4576
rect 5813 4573 5825 4576
rect 5859 4573 5871 4607
rect 6012 4604 6040 4635
rect 6178 4632 6184 4684
rect 6236 4632 6242 4684
rect 6822 4632 6828 4684
rect 6880 4632 6886 4684
rect 9030 4681 9036 4684
rect 7745 4675 7803 4681
rect 7745 4641 7757 4675
rect 7791 4672 7803 4675
rect 9008 4675 9036 4681
rect 7791 4644 8340 4672
rect 7791 4641 7803 4644
rect 7745 4635 7803 4641
rect 6840 4604 6868 4632
rect 7929 4607 7987 4613
rect 7929 4604 7941 4607
rect 6012 4576 6868 4604
rect 7852 4576 7941 4604
rect 5813 4567 5871 4573
rect 2133 4539 2191 4545
rect 2133 4505 2145 4539
rect 2179 4536 2191 4539
rect 3510 4536 3516 4548
rect 2179 4508 3516 4536
rect 2179 4505 2191 4508
rect 2133 4499 2191 4505
rect 3510 4496 3516 4508
rect 3568 4496 3574 4548
rect 4246 4496 4252 4548
rect 4304 4536 4310 4548
rect 4522 4536 4528 4548
rect 4304 4508 4528 4536
rect 4304 4496 4310 4508
rect 4522 4496 4528 4508
rect 4580 4536 4586 4548
rect 6178 4536 6184 4548
rect 4580 4508 6184 4536
rect 4580 4496 4586 4508
rect 6178 4496 6184 4508
rect 6236 4496 6242 4548
rect 4890 4428 4896 4480
rect 4948 4468 4954 4480
rect 7006 4468 7012 4480
rect 4948 4440 7012 4468
rect 4948 4428 4954 4440
rect 7006 4428 7012 4440
rect 7064 4468 7070 4480
rect 7852 4468 7880 4576
rect 7929 4573 7941 4576
rect 7975 4604 7987 4607
rect 8202 4604 8208 4616
rect 7975 4576 8208 4604
rect 7975 4573 7987 4576
rect 7929 4567 7987 4573
rect 8202 4564 8208 4576
rect 8260 4564 8266 4616
rect 7064 4440 7880 4468
rect 8312 4468 8340 4644
rect 9008 4641 9020 4675
rect 9008 4635 9036 4641
rect 9030 4632 9036 4635
rect 9088 4632 9094 4684
rect 9122 4632 9128 4684
rect 9180 4632 9186 4684
rect 9861 4675 9919 4681
rect 9861 4641 9873 4675
rect 9907 4672 9919 4675
rect 10137 4675 10195 4681
rect 10137 4672 10149 4675
rect 9907 4644 10149 4672
rect 9907 4641 9919 4644
rect 9861 4635 9919 4641
rect 10137 4641 10149 4644
rect 10183 4641 10195 4675
rect 10137 4635 10195 4641
rect 8662 4564 8668 4616
rect 8720 4604 8726 4616
rect 8849 4607 8907 4613
rect 8849 4604 8861 4607
rect 8720 4576 8861 4604
rect 8720 4564 8726 4576
rect 8849 4573 8861 4576
rect 8895 4573 8907 4607
rect 8849 4567 8907 4573
rect 9401 4607 9459 4613
rect 9401 4573 9413 4607
rect 9447 4604 9459 4607
rect 9950 4604 9956 4616
rect 9447 4576 9956 4604
rect 9447 4573 9459 4576
rect 9401 4567 9459 4573
rect 9950 4564 9956 4576
rect 10008 4564 10014 4616
rect 10045 4607 10103 4613
rect 10045 4573 10057 4607
rect 10091 4604 10103 4607
rect 10244 4604 10272 4712
rect 10594 4700 10600 4712
rect 10652 4700 10658 4752
rect 10321 4675 10379 4681
rect 10321 4641 10333 4675
rect 10367 4672 10379 4675
rect 11164 4672 11192 4780
rect 11238 4768 11244 4780
rect 11296 4768 11302 4820
rect 11514 4768 11520 4820
rect 11572 4808 11578 4820
rect 13817 4811 13875 4817
rect 13817 4808 13829 4811
rect 11572 4780 13829 4808
rect 11572 4768 11578 4780
rect 13817 4777 13829 4780
rect 13863 4808 13875 4811
rect 14182 4808 14188 4820
rect 13863 4780 14188 4808
rect 13863 4777 13875 4780
rect 13817 4771 13875 4777
rect 14182 4768 14188 4780
rect 14240 4768 14246 4820
rect 11422 4700 11428 4752
rect 11480 4740 11486 4752
rect 11480 4712 11928 4740
rect 11480 4700 11486 4712
rect 10367 4644 11192 4672
rect 10367 4641 10379 4644
rect 10321 4635 10379 4641
rect 11238 4632 11244 4684
rect 11296 4672 11302 4684
rect 11900 4681 11928 4712
rect 12066 4700 12072 4752
rect 12124 4740 12130 4752
rect 13265 4743 13323 4749
rect 13265 4740 13277 4743
rect 12124 4712 13277 4740
rect 12124 4700 12130 4712
rect 13265 4709 13277 4712
rect 13311 4709 13323 4743
rect 13265 4703 13323 4709
rect 11333 4675 11391 4681
rect 11333 4672 11345 4675
rect 11296 4644 11345 4672
rect 11296 4632 11302 4644
rect 11333 4641 11345 4644
rect 11379 4641 11391 4675
rect 11333 4635 11391 4641
rect 11885 4675 11943 4681
rect 11885 4641 11897 4675
rect 11931 4672 11943 4675
rect 12618 4672 12624 4684
rect 11931 4644 12624 4672
rect 11931 4641 11943 4644
rect 11885 4635 11943 4641
rect 12618 4632 12624 4644
rect 12676 4632 12682 4684
rect 12894 4632 12900 4684
rect 12952 4632 12958 4684
rect 13170 4632 13176 4684
rect 13228 4632 13234 4684
rect 14001 4675 14059 4681
rect 14001 4641 14013 4675
rect 14047 4672 14059 4675
rect 14366 4672 14372 4684
rect 14047 4644 14372 4672
rect 14047 4641 14059 4644
rect 14001 4635 14059 4641
rect 14366 4632 14372 4644
rect 14424 4632 14430 4684
rect 14642 4632 14648 4684
rect 14700 4672 14706 4684
rect 14921 4675 14979 4681
rect 14921 4672 14933 4675
rect 14700 4644 14933 4672
rect 14700 4632 14706 4644
rect 14921 4641 14933 4644
rect 14967 4641 14979 4675
rect 14921 4635 14979 4641
rect 10091 4576 10272 4604
rect 10505 4607 10563 4613
rect 10091 4573 10103 4576
rect 10045 4567 10103 4573
rect 10505 4573 10517 4607
rect 10551 4573 10563 4607
rect 10505 4567 10563 4573
rect 11425 4607 11483 4613
rect 11425 4573 11437 4607
rect 11471 4604 11483 4607
rect 11514 4604 11520 4616
rect 11471 4576 11520 4604
rect 11471 4573 11483 4576
rect 11425 4567 11483 4573
rect 9490 4496 9496 4548
rect 9548 4536 9554 4548
rect 10520 4536 10548 4567
rect 11514 4564 11520 4576
rect 11572 4564 11578 4616
rect 11609 4607 11667 4613
rect 11609 4573 11621 4607
rect 11655 4604 11667 4607
rect 12158 4604 12164 4616
rect 11655 4576 12164 4604
rect 11655 4573 11667 4576
rect 11609 4567 11667 4573
rect 12158 4564 12164 4576
rect 12216 4564 12222 4616
rect 12250 4564 12256 4616
rect 12308 4604 12314 4616
rect 12437 4607 12495 4613
rect 12437 4604 12449 4607
rect 12308 4576 12449 4604
rect 12308 4564 12314 4576
rect 12437 4573 12449 4576
rect 12483 4604 12495 4607
rect 12912 4604 12940 4632
rect 12483 4576 12940 4604
rect 12483 4573 12495 4576
rect 12437 4567 12495 4573
rect 13078 4564 13084 4616
rect 13136 4564 13142 4616
rect 13357 4607 13415 4613
rect 13357 4573 13369 4607
rect 13403 4573 13415 4607
rect 13357 4567 13415 4573
rect 9548 4508 10548 4536
rect 9548 4496 9554 4508
rect 10778 4496 10784 4548
rect 10836 4536 10842 4548
rect 13096 4536 13124 4564
rect 10836 4508 13124 4536
rect 10836 4496 10842 4508
rect 10042 4468 10048 4480
rect 8312 4440 10048 4468
rect 7064 4428 7070 4440
rect 10042 4428 10048 4440
rect 10100 4428 10106 4480
rect 10870 4428 10876 4480
rect 10928 4468 10934 4480
rect 12066 4468 12072 4480
rect 10928 4440 12072 4468
rect 10928 4428 10934 4440
rect 12066 4428 12072 4440
rect 12124 4428 12130 4480
rect 12802 4428 12808 4480
rect 12860 4428 12866 4480
rect 13078 4428 13084 4480
rect 13136 4468 13142 4480
rect 13372 4468 13400 4567
rect 14458 4564 14464 4616
rect 14516 4564 14522 4616
rect 13136 4440 13400 4468
rect 13136 4428 13142 4440
rect 552 4378 15364 4400
rect 552 4326 2249 4378
rect 2301 4326 2313 4378
rect 2365 4326 2377 4378
rect 2429 4326 2441 4378
rect 2493 4326 2505 4378
rect 2557 4326 5951 4378
rect 6003 4326 6015 4378
rect 6067 4326 6079 4378
rect 6131 4326 6143 4378
rect 6195 4326 6207 4378
rect 6259 4326 9653 4378
rect 9705 4326 9717 4378
rect 9769 4326 9781 4378
rect 9833 4326 9845 4378
rect 9897 4326 9909 4378
rect 9961 4326 13355 4378
rect 13407 4326 13419 4378
rect 13471 4326 13483 4378
rect 13535 4326 13547 4378
rect 13599 4326 13611 4378
rect 13663 4326 15364 4378
rect 552 4304 15364 4326
rect 3697 4267 3755 4273
rect 3697 4233 3709 4267
rect 3743 4264 3755 4267
rect 4338 4264 4344 4276
rect 3743 4236 4344 4264
rect 3743 4233 3755 4236
rect 3697 4227 3755 4233
rect 4338 4224 4344 4236
rect 4396 4224 4402 4276
rect 9398 4264 9404 4276
rect 8588 4236 9404 4264
rect 2501 4199 2559 4205
rect 2501 4165 2513 4199
rect 2547 4196 2559 4199
rect 6730 4196 6736 4208
rect 2547 4168 3372 4196
rect 2547 4165 2559 4168
rect 2501 4159 2559 4165
rect 2225 4131 2283 4137
rect 2225 4097 2237 4131
rect 2271 4128 2283 4131
rect 2682 4128 2688 4140
rect 2271 4100 2688 4128
rect 2271 4097 2283 4100
rect 2225 4091 2283 4097
rect 2682 4088 2688 4100
rect 2740 4088 2746 4140
rect 3344 4137 3372 4168
rect 6012 4168 6736 4196
rect 3329 4131 3387 4137
rect 3329 4097 3341 4131
rect 3375 4097 3387 4131
rect 3329 4091 3387 4097
rect 4246 4088 4252 4140
rect 4304 4088 4310 4140
rect 4430 4088 4436 4140
rect 4488 4128 4494 4140
rect 6012 4137 6040 4168
rect 6730 4156 6736 4168
rect 6788 4196 6794 4208
rect 6917 4199 6975 4205
rect 6917 4196 6929 4199
rect 6788 4168 6929 4196
rect 6788 4156 6794 4168
rect 6917 4165 6929 4168
rect 6963 4196 6975 4199
rect 7006 4196 7012 4208
rect 6963 4168 7012 4196
rect 6963 4165 6975 4168
rect 6917 4159 6975 4165
rect 7006 4156 7012 4168
rect 7064 4156 7070 4208
rect 8588 4137 8616 4236
rect 9398 4224 9404 4236
rect 9456 4264 9462 4276
rect 10134 4264 10140 4276
rect 9456 4236 10140 4264
rect 9456 4224 9462 4236
rect 10134 4224 10140 4236
rect 10192 4224 10198 4276
rect 10597 4267 10655 4273
rect 10597 4233 10609 4267
rect 10643 4264 10655 4267
rect 10870 4264 10876 4276
rect 10643 4236 10876 4264
rect 10643 4233 10655 4236
rect 10597 4227 10655 4233
rect 10870 4224 10876 4236
rect 10928 4224 10934 4276
rect 11514 4224 11520 4276
rect 11572 4264 11578 4276
rect 11701 4267 11759 4273
rect 11701 4264 11713 4267
rect 11572 4236 11713 4264
rect 11572 4224 11578 4236
rect 11701 4233 11713 4236
rect 11747 4233 11759 4267
rect 11701 4227 11759 4233
rect 9122 4156 9128 4208
rect 9180 4156 9186 4208
rect 12268 4168 13032 4196
rect 4709 4131 4767 4137
rect 4709 4128 4721 4131
rect 4488 4100 4721 4128
rect 4488 4088 4494 4100
rect 4709 4097 4721 4100
rect 4755 4097 4767 4131
rect 4709 4091 4767 4097
rect 5997 4131 6055 4137
rect 5997 4097 6009 4131
rect 6043 4097 6055 4131
rect 6411 4131 6469 4137
rect 6411 4128 6423 4131
rect 5997 4091 6055 4097
rect 6104 4100 6423 4128
rect 2133 4063 2191 4069
rect 2133 4029 2145 4063
rect 2179 4060 2191 4063
rect 2590 4060 2596 4072
rect 2179 4032 2596 4060
rect 2179 4029 2191 4032
rect 2133 4023 2191 4029
rect 2590 4020 2596 4032
rect 2648 4020 2654 4072
rect 3234 4020 3240 4072
rect 3292 4060 3298 4072
rect 3421 4063 3479 4069
rect 3421 4060 3433 4063
rect 3292 4032 3433 4060
rect 3292 4020 3298 4032
rect 3421 4029 3433 4032
rect 3467 4060 3479 4063
rect 3970 4060 3976 4072
rect 3467 4032 3976 4060
rect 3467 4029 3479 4032
rect 3421 4023 3479 4029
rect 3970 4020 3976 4032
rect 4028 4020 4034 4072
rect 4062 4020 4068 4072
rect 4120 4020 4126 4072
rect 5718 4060 5724 4072
rect 5000 4032 5724 4060
rect 5000 4001 5028 4032
rect 5718 4020 5724 4032
rect 5776 4060 5782 4072
rect 6104 4060 6132 4100
rect 6411 4097 6423 4100
rect 6457 4097 6469 4131
rect 7310 4131 7368 4137
rect 7310 4128 7322 4131
rect 6411 4091 6469 4097
rect 6656 4100 7322 4128
rect 6656 4072 6684 4100
rect 7310 4097 7322 4100
rect 7356 4097 7368 4131
rect 7310 4091 7368 4097
rect 8573 4131 8631 4137
rect 8573 4097 8585 4131
rect 8619 4097 8631 4131
rect 8573 4091 8631 4097
rect 8665 4131 8723 4137
rect 8665 4097 8677 4131
rect 8711 4128 8723 4131
rect 8754 4128 8760 4140
rect 8711 4100 8760 4128
rect 8711 4097 8723 4100
rect 8665 4091 8723 4097
rect 8754 4088 8760 4100
rect 8812 4088 8818 4140
rect 8956 4100 9674 4128
rect 5776 4032 6132 4060
rect 5776 4020 5782 4032
rect 6178 4020 6184 4072
rect 6236 4060 6242 4072
rect 6273 4063 6331 4069
rect 6273 4060 6285 4063
rect 6236 4032 6285 4060
rect 6236 4020 6242 4032
rect 6273 4029 6285 4032
rect 6319 4029 6331 4063
rect 6273 4023 6331 4029
rect 6638 4020 6644 4072
rect 6696 4020 6702 4072
rect 7190 4020 7196 4072
rect 7248 4020 7254 4072
rect 7466 4020 7472 4072
rect 7524 4020 7530 4072
rect 8113 4063 8171 4069
rect 8113 4029 8125 4063
rect 8159 4060 8171 4063
rect 8956 4060 8984 4100
rect 8159 4032 8984 4060
rect 8159 4029 8171 4032
rect 8113 4023 8171 4029
rect 9122 4020 9128 4072
rect 9180 4060 9186 4072
rect 9401 4063 9459 4069
rect 9401 4060 9413 4063
rect 9180 4032 9413 4060
rect 9180 4020 9186 4032
rect 9401 4029 9413 4032
rect 9447 4029 9459 4063
rect 9646 4060 9674 4100
rect 10042 4088 10048 4140
rect 10100 4128 10106 4140
rect 10873 4131 10931 4137
rect 10873 4128 10885 4131
rect 10100 4100 10885 4128
rect 10100 4088 10106 4100
rect 10873 4097 10885 4100
rect 10919 4128 10931 4131
rect 12158 4128 12164 4140
rect 10919 4100 12164 4128
rect 10919 4097 10931 4100
rect 10873 4091 10931 4097
rect 12158 4088 12164 4100
rect 12216 4088 12222 4140
rect 10137 4063 10195 4069
rect 10137 4060 10149 4063
rect 9646 4032 10149 4060
rect 9401 4023 9459 4029
rect 10137 4029 10149 4032
rect 10183 4029 10195 4063
rect 10137 4023 10195 4029
rect 10226 4020 10232 4072
rect 10284 4020 10290 4072
rect 11054 4020 11060 4072
rect 11112 4020 11118 4072
rect 12268 4060 12296 4168
rect 12345 4131 12403 4137
rect 12345 4097 12357 4131
rect 12391 4128 12403 4131
rect 12526 4128 12532 4140
rect 12391 4100 12532 4128
rect 12391 4097 12403 4100
rect 12345 4091 12403 4097
rect 12526 4088 12532 4100
rect 12584 4128 12590 4140
rect 12710 4128 12716 4140
rect 12584 4100 12716 4128
rect 12584 4088 12590 4100
rect 12710 4088 12716 4100
rect 12768 4088 12774 4140
rect 12802 4088 12808 4140
rect 12860 4088 12866 4140
rect 13004 4137 13032 4168
rect 12989 4131 13047 4137
rect 12989 4097 13001 4131
rect 13035 4097 13047 4131
rect 12989 4091 13047 4097
rect 13078 4088 13084 4140
rect 13136 4088 13142 4140
rect 14090 4128 14096 4140
rect 13188 4100 14096 4128
rect 11440 4032 12296 4060
rect 12820 4060 12848 4088
rect 12897 4063 12955 4069
rect 12897 4060 12909 4063
rect 12820 4032 12909 4060
rect 4985 3995 5043 4001
rect 4985 3992 4997 3995
rect 3436 3964 4997 3992
rect 3436 3936 3464 3964
rect 4985 3961 4997 3964
rect 5031 3961 5043 3995
rect 8757 3995 8815 4001
rect 8757 3992 8769 3995
rect 4985 3955 5043 3961
rect 7944 3964 8769 3992
rect 3418 3884 3424 3936
rect 3476 3884 3482 3936
rect 3878 3884 3884 3936
rect 3936 3884 3942 3936
rect 4890 3884 4896 3936
rect 4948 3884 4954 3936
rect 5350 3884 5356 3936
rect 5408 3884 5414 3936
rect 5442 3884 5448 3936
rect 5500 3884 5506 3936
rect 5810 3884 5816 3936
rect 5868 3884 5874 3936
rect 5905 3927 5963 3933
rect 5905 3893 5917 3927
rect 5951 3924 5963 3927
rect 7190 3924 7196 3936
rect 5951 3896 7196 3924
rect 5951 3893 5963 3896
rect 5905 3887 5963 3893
rect 7190 3884 7196 3896
rect 7248 3884 7254 3936
rect 7466 3884 7472 3936
rect 7524 3924 7530 3936
rect 7944 3924 7972 3964
rect 8757 3961 8769 3964
rect 8803 3961 8815 3995
rect 11072 3992 11100 4020
rect 8757 3955 8815 3961
rect 9646 3964 11100 3992
rect 7524 3896 7972 3924
rect 7524 3884 7530 3896
rect 9214 3884 9220 3936
rect 9272 3884 9278 3936
rect 9398 3884 9404 3936
rect 9456 3924 9462 3936
rect 9646 3924 9674 3964
rect 9456 3896 9674 3924
rect 9456 3884 9462 3896
rect 9766 3884 9772 3936
rect 9824 3924 9830 3936
rect 10962 3924 10968 3936
rect 9824 3896 10968 3924
rect 9824 3884 9830 3896
rect 10962 3884 10968 3896
rect 11020 3884 11026 3936
rect 11054 3884 11060 3936
rect 11112 3884 11118 3936
rect 11440 3933 11468 4032
rect 12897 4029 12909 4032
rect 12943 4029 12955 4063
rect 12897 4023 12955 4029
rect 11882 3952 11888 4004
rect 11940 3992 11946 4004
rect 12069 3995 12127 4001
rect 12069 3992 12081 3995
rect 11940 3964 12081 3992
rect 11940 3952 11946 3964
rect 12069 3961 12081 3964
rect 12115 3992 12127 3995
rect 13188 3992 13216 4100
rect 14090 4088 14096 4100
rect 14148 4088 14154 4140
rect 14642 4088 14648 4140
rect 14700 4128 14706 4140
rect 14737 4131 14795 4137
rect 14737 4128 14749 4131
rect 14700 4100 14749 4128
rect 14700 4088 14706 4100
rect 14737 4097 14749 4100
rect 14783 4097 14795 4131
rect 14737 4091 14795 4097
rect 13906 4020 13912 4072
rect 13964 4020 13970 4072
rect 13998 4020 14004 4072
rect 14056 4020 14062 4072
rect 15013 4063 15071 4069
rect 15013 4029 15025 4063
rect 15059 4060 15071 4063
rect 15102 4060 15108 4072
rect 15059 4032 15108 4060
rect 15059 4029 15071 4032
rect 15013 4023 15071 4029
rect 15102 4020 15108 4032
rect 15160 4020 15166 4072
rect 12115 3964 13216 3992
rect 12115 3961 12127 3964
rect 12069 3955 12127 3961
rect 13354 3952 13360 4004
rect 13412 3992 13418 4004
rect 14016 3992 14044 4020
rect 13412 3964 13952 3992
rect 14016 3964 14596 3992
rect 13412 3952 13418 3964
rect 11425 3927 11483 3933
rect 11425 3893 11437 3927
rect 11471 3893 11483 3927
rect 11425 3887 11483 3893
rect 12158 3884 12164 3936
rect 12216 3884 12222 3936
rect 12250 3884 12256 3936
rect 12308 3924 12314 3936
rect 12529 3927 12587 3933
rect 12529 3924 12541 3927
rect 12308 3896 12541 3924
rect 12308 3884 12314 3896
rect 12529 3893 12541 3896
rect 12575 3893 12587 3927
rect 12529 3887 12587 3893
rect 13170 3884 13176 3936
rect 13228 3924 13234 3936
rect 13541 3927 13599 3933
rect 13541 3924 13553 3927
rect 13228 3896 13553 3924
rect 13228 3884 13234 3896
rect 13541 3893 13553 3896
rect 13587 3893 13599 3927
rect 13924 3924 13952 3964
rect 14568 3936 14596 3964
rect 14001 3927 14059 3933
rect 14001 3924 14013 3927
rect 13924 3896 14013 3924
rect 13541 3887 13599 3893
rect 14001 3893 14013 3896
rect 14047 3893 14059 3927
rect 14001 3887 14059 3893
rect 14550 3884 14556 3936
rect 14608 3884 14614 3936
rect 14826 3884 14832 3936
rect 14884 3924 14890 3936
rect 15102 3924 15108 3936
rect 14884 3896 15108 3924
rect 14884 3884 14890 3896
rect 15102 3884 15108 3896
rect 15160 3884 15166 3936
rect 552 3834 15520 3856
rect 552 3782 4100 3834
rect 4152 3782 4164 3834
rect 4216 3782 4228 3834
rect 4280 3782 4292 3834
rect 4344 3782 4356 3834
rect 4408 3782 7802 3834
rect 7854 3782 7866 3834
rect 7918 3782 7930 3834
rect 7982 3782 7994 3834
rect 8046 3782 8058 3834
rect 8110 3782 11504 3834
rect 11556 3782 11568 3834
rect 11620 3782 11632 3834
rect 11684 3782 11696 3834
rect 11748 3782 11760 3834
rect 11812 3782 15206 3834
rect 15258 3782 15270 3834
rect 15322 3782 15334 3834
rect 15386 3782 15398 3834
rect 15450 3782 15462 3834
rect 15514 3782 15520 3834
rect 552 3760 15520 3782
rect 3421 3723 3479 3729
rect 3421 3689 3433 3723
rect 3467 3720 3479 3723
rect 3602 3720 3608 3732
rect 3467 3692 3608 3720
rect 3467 3689 3479 3692
rect 3421 3683 3479 3689
rect 3602 3680 3608 3692
rect 3660 3680 3666 3732
rect 5810 3720 5816 3732
rect 3804 3692 5816 3720
rect 1118 3544 1124 3596
rect 1176 3584 1182 3596
rect 3804 3593 3832 3692
rect 5810 3680 5816 3692
rect 5868 3720 5874 3732
rect 6638 3720 6644 3732
rect 5868 3692 6644 3720
rect 5868 3680 5874 3692
rect 6638 3680 6644 3692
rect 6696 3680 6702 3732
rect 8846 3680 8852 3732
rect 8904 3680 8910 3732
rect 9858 3680 9864 3732
rect 9916 3680 9922 3732
rect 10042 3680 10048 3732
rect 10100 3720 10106 3732
rect 10229 3723 10287 3729
rect 10229 3720 10241 3723
rect 10100 3692 10241 3720
rect 10100 3680 10106 3692
rect 10229 3689 10241 3692
rect 10275 3689 10287 3723
rect 10229 3683 10287 3689
rect 11146 3680 11152 3732
rect 11204 3720 11210 3732
rect 11790 3720 11796 3732
rect 11204 3692 11796 3720
rect 11204 3680 11210 3692
rect 11790 3680 11796 3692
rect 11848 3680 11854 3732
rect 12986 3680 12992 3732
rect 13044 3720 13050 3732
rect 13044 3692 13400 3720
rect 13044 3680 13050 3692
rect 5074 3612 5080 3664
rect 5132 3652 5138 3664
rect 5132 3624 5948 3652
rect 5132 3612 5138 3624
rect 3789 3587 3847 3593
rect 3789 3584 3801 3587
rect 1176 3556 3801 3584
rect 1176 3544 1182 3556
rect 3789 3553 3801 3556
rect 3835 3553 3847 3587
rect 3789 3547 3847 3553
rect 3970 3544 3976 3596
rect 4028 3584 4034 3596
rect 4985 3587 5043 3593
rect 4985 3584 4997 3587
rect 4028 3556 4997 3584
rect 4028 3544 4034 3556
rect 4985 3553 4997 3556
rect 5031 3553 5043 3587
rect 4985 3547 5043 3553
rect 5169 3587 5227 3593
rect 5169 3553 5181 3587
rect 5215 3584 5227 3587
rect 5350 3584 5356 3596
rect 5215 3556 5356 3584
rect 5215 3553 5227 3556
rect 5169 3547 5227 3553
rect 3050 3476 3056 3528
rect 3108 3516 3114 3528
rect 3881 3519 3939 3525
rect 3881 3516 3893 3519
rect 3108 3488 3893 3516
rect 3108 3476 3114 3488
rect 3881 3485 3893 3488
rect 3927 3485 3939 3519
rect 3881 3479 3939 3485
rect 4065 3519 4123 3525
rect 4065 3485 4077 3519
rect 4111 3516 4123 3519
rect 4338 3516 4344 3528
rect 4111 3488 4344 3516
rect 4111 3485 4123 3488
rect 4065 3479 4123 3485
rect 4338 3476 4344 3488
rect 4396 3476 4402 3528
rect 5000 3516 5028 3547
rect 5350 3544 5356 3556
rect 5408 3544 5414 3596
rect 5442 3544 5448 3596
rect 5500 3584 5506 3596
rect 5813 3587 5871 3593
rect 5813 3584 5825 3587
rect 5500 3556 5825 3584
rect 5500 3544 5506 3556
rect 5813 3553 5825 3556
rect 5859 3553 5871 3587
rect 5920 3584 5948 3624
rect 6178 3612 6184 3664
rect 6236 3652 6242 3664
rect 6730 3652 6736 3664
rect 6236 3624 6736 3652
rect 6236 3612 6242 3624
rect 6730 3612 6736 3624
rect 6788 3612 6794 3664
rect 7374 3612 7380 3664
rect 7432 3652 7438 3664
rect 9674 3652 9680 3664
rect 7432 3624 9680 3652
rect 7432 3612 7438 3624
rect 9674 3612 9680 3624
rect 9732 3612 9738 3664
rect 9876 3652 9904 3680
rect 9784 3624 9904 3652
rect 8754 3584 8760 3596
rect 5920 3556 8760 3584
rect 5813 3547 5871 3553
rect 8754 3544 8760 3556
rect 8812 3544 8818 3596
rect 9582 3544 9588 3596
rect 9640 3544 9646 3596
rect 9784 3593 9812 3624
rect 12526 3612 12532 3664
rect 12584 3652 12590 3664
rect 13078 3652 13084 3664
rect 12584 3624 13084 3652
rect 12584 3612 12590 3624
rect 13078 3612 13084 3624
rect 13136 3612 13142 3664
rect 9769 3587 9827 3593
rect 9769 3553 9781 3587
rect 9815 3553 9827 3587
rect 9769 3547 9827 3553
rect 11793 3587 11851 3593
rect 11793 3553 11805 3587
rect 11839 3584 11851 3587
rect 11882 3584 11888 3596
rect 11839 3556 11888 3584
rect 11839 3553 11851 3556
rect 11793 3547 11851 3553
rect 11882 3544 11888 3556
rect 11940 3544 11946 3596
rect 11974 3544 11980 3596
rect 12032 3544 12038 3596
rect 13170 3544 13176 3596
rect 13228 3544 13234 3596
rect 13372 3593 13400 3692
rect 13906 3680 13912 3732
rect 13964 3720 13970 3732
rect 15013 3723 15071 3729
rect 15013 3720 15025 3723
rect 13964 3692 15025 3720
rect 13964 3680 13970 3692
rect 15013 3689 15025 3692
rect 15059 3689 15071 3723
rect 15013 3683 15071 3689
rect 13357 3587 13415 3593
rect 13357 3553 13369 3587
rect 13403 3553 13415 3587
rect 13357 3547 13415 3553
rect 14090 3544 14096 3596
rect 14148 3544 14154 3596
rect 5534 3516 5540 3528
rect 5000 3488 5540 3516
rect 5534 3476 5540 3488
rect 5592 3476 5598 3528
rect 9033 3519 9091 3525
rect 9033 3485 9045 3519
rect 9079 3516 9091 3519
rect 9079 3488 9904 3516
rect 9079 3485 9091 3488
rect 9033 3479 9091 3485
rect 5353 3451 5411 3457
rect 5353 3417 5365 3451
rect 5399 3448 5411 3451
rect 9766 3448 9772 3460
rect 5399 3420 9772 3448
rect 5399 3417 5411 3420
rect 5353 3411 5411 3417
rect 9766 3408 9772 3420
rect 9824 3408 9830 3460
rect 9876 3448 9904 3488
rect 11238 3476 11244 3528
rect 11296 3516 11302 3528
rect 14210 3519 14268 3525
rect 14210 3516 14222 3519
rect 11296 3488 14222 3516
rect 11296 3476 11302 3488
rect 14210 3485 14222 3488
rect 14256 3485 14268 3519
rect 14210 3479 14268 3485
rect 14369 3519 14427 3525
rect 14369 3485 14381 3519
rect 14415 3516 14427 3519
rect 14415 3488 14780 3516
rect 14415 3485 14427 3488
rect 14369 3479 14427 3485
rect 11146 3448 11152 3460
rect 9876 3420 11152 3448
rect 11146 3408 11152 3420
rect 11204 3408 11210 3460
rect 12158 3408 12164 3460
rect 12216 3408 12222 3460
rect 12250 3408 12256 3460
rect 12308 3448 12314 3460
rect 13817 3451 13875 3457
rect 13817 3448 13829 3451
rect 12308 3420 13829 3448
rect 12308 3408 12314 3420
rect 13817 3417 13829 3420
rect 13863 3417 13875 3451
rect 13817 3411 13875 3417
rect 3142 3340 3148 3392
rect 3200 3380 3206 3392
rect 4801 3383 4859 3389
rect 4801 3380 4813 3383
rect 3200 3352 4813 3380
rect 3200 3340 3206 3352
rect 4801 3349 4813 3352
rect 4847 3349 4859 3383
rect 4801 3343 4859 3349
rect 5810 3340 5816 3392
rect 5868 3380 5874 3392
rect 5997 3383 6055 3389
rect 5997 3380 6009 3383
rect 5868 3352 6009 3380
rect 5868 3340 5874 3352
rect 5997 3349 6009 3352
rect 6043 3349 6055 3383
rect 5997 3343 6055 3349
rect 8386 3340 8392 3392
rect 8444 3340 8450 3392
rect 8478 3340 8484 3392
rect 8536 3380 8542 3392
rect 9674 3380 9680 3392
rect 8536 3352 9680 3380
rect 8536 3340 8542 3352
rect 9674 3340 9680 3352
rect 9732 3340 9738 3392
rect 9861 3383 9919 3389
rect 9861 3349 9873 3383
rect 9907 3380 9919 3383
rect 10962 3380 10968 3392
rect 9907 3352 10968 3380
rect 9907 3349 9919 3352
rect 9861 3343 9919 3349
rect 10962 3340 10968 3352
rect 11020 3340 11026 3392
rect 12069 3383 12127 3389
rect 12069 3349 12081 3383
rect 12115 3380 12127 3383
rect 12176 3380 12204 3408
rect 12115 3352 12204 3380
rect 12115 3349 12127 3352
rect 12069 3343 12127 3349
rect 13170 3340 13176 3392
rect 13228 3380 13234 3392
rect 13354 3380 13360 3392
rect 13228 3352 13360 3380
rect 13228 3340 13234 3352
rect 13354 3340 13360 3352
rect 13412 3340 13418 3392
rect 14182 3340 14188 3392
rect 14240 3380 14246 3392
rect 14752 3380 14780 3488
rect 14240 3352 14780 3380
rect 14240 3340 14246 3352
rect 552 3290 15364 3312
rect 552 3238 2249 3290
rect 2301 3238 2313 3290
rect 2365 3238 2377 3290
rect 2429 3238 2441 3290
rect 2493 3238 2505 3290
rect 2557 3238 5951 3290
rect 6003 3238 6015 3290
rect 6067 3238 6079 3290
rect 6131 3238 6143 3290
rect 6195 3238 6207 3290
rect 6259 3238 9653 3290
rect 9705 3238 9717 3290
rect 9769 3238 9781 3290
rect 9833 3238 9845 3290
rect 9897 3238 9909 3290
rect 9961 3238 13355 3290
rect 13407 3238 13419 3290
rect 13471 3238 13483 3290
rect 13535 3238 13547 3290
rect 13599 3238 13611 3290
rect 13663 3238 15364 3290
rect 552 3216 15364 3238
rect 4982 3136 4988 3188
rect 5040 3136 5046 3188
rect 6365 3179 6423 3185
rect 6365 3145 6377 3179
rect 6411 3176 6423 3179
rect 7374 3176 7380 3188
rect 6411 3148 7380 3176
rect 6411 3145 6423 3148
rect 6365 3139 6423 3145
rect 7374 3136 7380 3148
rect 7432 3136 7438 3188
rect 8846 3136 8852 3188
rect 8904 3176 8910 3188
rect 8904 3148 9352 3176
rect 8904 3136 8910 3148
rect 7006 3068 7012 3120
rect 7064 3108 7070 3120
rect 7064 3080 7144 3108
rect 7064 3068 7070 3080
rect 4338 3000 4344 3052
rect 4396 3000 4402 3052
rect 5718 3000 5724 3052
rect 5776 3040 5782 3052
rect 5776 3012 6224 3040
rect 5776 3000 5782 3012
rect 3234 2932 3240 2984
rect 3292 2972 3298 2984
rect 5810 2972 5816 2984
rect 3292 2944 5816 2972
rect 3292 2932 3298 2944
rect 5810 2932 5816 2944
rect 5868 2932 5874 2984
rect 5902 2932 5908 2984
rect 5960 2932 5966 2984
rect 6089 2975 6147 2981
rect 6089 2941 6101 2975
rect 6135 2941 6147 2975
rect 6196 2972 6224 3012
rect 6730 3000 6736 3052
rect 6788 3040 6794 3052
rect 7116 3049 7144 3080
rect 7101 3043 7159 3049
rect 6788 3012 7052 3040
rect 6788 3000 6794 3012
rect 7024 2981 7052 3012
rect 7101 3009 7113 3043
rect 7147 3009 7159 3043
rect 7101 3003 7159 3009
rect 8478 3000 8484 3052
rect 8536 3000 8542 3052
rect 8938 3000 8944 3052
rect 8996 3040 9002 3052
rect 9217 3043 9275 3049
rect 9217 3040 9229 3043
rect 8996 3012 9229 3040
rect 8996 3000 9002 3012
rect 9217 3009 9229 3012
rect 9263 3009 9275 3043
rect 9324 3040 9352 3148
rect 10226 3136 10232 3188
rect 10284 3176 10290 3188
rect 10413 3179 10471 3185
rect 10413 3176 10425 3179
rect 10284 3148 10425 3176
rect 10284 3136 10290 3148
rect 10413 3145 10425 3148
rect 10459 3145 10471 3179
rect 10413 3139 10471 3145
rect 11333 3179 11391 3185
rect 11333 3145 11345 3179
rect 11379 3176 11391 3179
rect 11974 3176 11980 3188
rect 11379 3148 11980 3176
rect 11379 3145 11391 3148
rect 11333 3139 11391 3145
rect 11974 3136 11980 3148
rect 12032 3136 12038 3188
rect 12894 3136 12900 3188
rect 12952 3176 12958 3188
rect 13541 3179 13599 3185
rect 13541 3176 13553 3179
rect 12952 3148 13553 3176
rect 12952 3136 12958 3148
rect 13541 3145 13553 3148
rect 13587 3145 13599 3179
rect 13541 3139 13599 3145
rect 11054 3108 11060 3120
rect 10796 3080 11060 3108
rect 9324 3012 9536 3040
rect 9217 3003 9275 3009
rect 6917 2975 6975 2981
rect 6917 2972 6929 2975
rect 6196 2944 6929 2972
rect 6089 2935 6147 2941
rect 6917 2941 6929 2944
rect 6963 2941 6975 2975
rect 6917 2935 6975 2941
rect 7009 2975 7067 2981
rect 7009 2941 7021 2975
rect 7055 2972 7067 2975
rect 8496 2972 8524 3000
rect 7055 2944 8524 2972
rect 8573 2975 8631 2981
rect 7055 2941 7067 2944
rect 7009 2935 7067 2941
rect 8573 2941 8585 2975
rect 8619 2941 8631 2975
rect 8573 2935 8631 2941
rect 5074 2904 5080 2916
rect 4632 2876 5080 2904
rect 3786 2796 3792 2848
rect 3844 2836 3850 2848
rect 4632 2845 4660 2876
rect 5074 2864 5080 2876
rect 5132 2864 5138 2916
rect 6104 2904 6132 2935
rect 7558 2904 7564 2916
rect 6104 2876 7564 2904
rect 7558 2864 7564 2876
rect 7616 2904 7622 2916
rect 8478 2904 8484 2916
rect 7616 2876 8484 2904
rect 7616 2864 7622 2876
rect 8478 2864 8484 2876
rect 8536 2864 8542 2916
rect 4525 2839 4583 2845
rect 4525 2836 4537 2839
rect 3844 2808 4537 2836
rect 3844 2796 3850 2808
rect 4525 2805 4537 2808
rect 4571 2805 4583 2839
rect 4525 2799 4583 2805
rect 4617 2839 4675 2845
rect 4617 2805 4629 2839
rect 4663 2805 4675 2839
rect 4617 2799 4675 2805
rect 6546 2796 6552 2848
rect 6604 2796 6610 2848
rect 8588 2836 8616 2935
rect 8754 2932 8760 2984
rect 8812 2932 8818 2984
rect 9508 2981 9536 3012
rect 9582 3000 9588 3052
rect 9640 3049 9646 3052
rect 10796 3049 10824 3080
rect 11054 3068 11060 3080
rect 11112 3068 11118 3120
rect 13170 3068 13176 3120
rect 13228 3108 13234 3120
rect 13357 3111 13415 3117
rect 13357 3108 13369 3111
rect 13228 3080 13369 3108
rect 13228 3068 13234 3080
rect 13357 3077 13369 3080
rect 13403 3077 13415 3111
rect 14369 3111 14427 3117
rect 14369 3108 14381 3111
rect 13357 3071 13415 3077
rect 14016 3080 14381 3108
rect 9640 3043 9668 3049
rect 9656 3009 9668 3043
rect 10781 3043 10839 3049
rect 10781 3040 10793 3043
rect 9640 3003 9668 3009
rect 9784 3012 10793 3040
rect 9640 3000 9646 3003
rect 9784 2984 9812 3012
rect 10781 3009 10793 3012
rect 10827 3009 10839 3043
rect 10781 3003 10839 3009
rect 11330 3000 11336 3052
rect 11388 3040 11394 3052
rect 11701 3043 11759 3049
rect 11701 3040 11713 3043
rect 11388 3012 11713 3040
rect 11388 3000 11394 3012
rect 11701 3009 11713 3012
rect 11747 3009 11759 3043
rect 11701 3003 11759 3009
rect 11790 3000 11796 3052
rect 11848 3040 11854 3052
rect 12161 3043 12219 3049
rect 12161 3040 12173 3043
rect 11848 3012 12173 3040
rect 11848 3000 11854 3012
rect 12161 3009 12173 3012
rect 12207 3040 12219 3043
rect 12250 3040 12256 3052
rect 12207 3012 12256 3040
rect 12207 3009 12219 3012
rect 12161 3003 12219 3009
rect 12250 3000 12256 3012
rect 12308 3000 12314 3052
rect 12434 3000 12440 3052
rect 12492 3040 12498 3052
rect 14016 3040 14044 3080
rect 14369 3077 14381 3080
rect 14415 3077 14427 3111
rect 14369 3071 14427 3077
rect 14642 3068 14648 3120
rect 14700 3068 14706 3120
rect 12492 3012 14044 3040
rect 12492 3000 12498 3012
rect 14090 3000 14096 3052
rect 14148 3000 14154 3052
rect 15562 3000 15568 3052
rect 15620 3000 15626 3052
rect 9493 2975 9551 2981
rect 9493 2941 9505 2975
rect 9539 2941 9551 2975
rect 9493 2935 9551 2941
rect 9766 2932 9772 2984
rect 9824 2932 9830 2984
rect 10870 2932 10876 2984
rect 10928 2932 10934 2984
rect 10962 2932 10968 2984
rect 11020 2972 11026 2984
rect 11057 2975 11115 2981
rect 11057 2972 11069 2975
rect 11020 2944 11069 2972
rect 11020 2932 11026 2944
rect 11057 2941 11069 2944
rect 11103 2941 11115 2975
rect 11057 2935 11115 2941
rect 11517 2975 11575 2981
rect 11517 2941 11529 2975
rect 11563 2941 11575 2975
rect 11517 2935 11575 2941
rect 10226 2836 10232 2848
rect 8588 2808 10232 2836
rect 10226 2796 10232 2808
rect 10284 2836 10290 2848
rect 10778 2836 10784 2848
rect 10284 2808 10784 2836
rect 10284 2796 10290 2808
rect 10778 2796 10784 2808
rect 10836 2796 10842 2848
rect 11532 2836 11560 2935
rect 12526 2932 12532 2984
rect 12584 2981 12590 2984
rect 12584 2975 12612 2981
rect 12600 2941 12612 2975
rect 12584 2935 12612 2941
rect 12584 2932 12590 2935
rect 12710 2932 12716 2984
rect 12768 2932 12774 2984
rect 14001 2975 14059 2981
rect 14001 2972 14013 2975
rect 13280 2944 14013 2972
rect 12250 2836 12256 2848
rect 11532 2808 12256 2836
rect 12250 2796 12256 2808
rect 12308 2796 12314 2848
rect 12710 2796 12716 2848
rect 12768 2836 12774 2848
rect 13280 2836 13308 2944
rect 14001 2941 14013 2944
rect 14047 2941 14059 2975
rect 14001 2935 14059 2941
rect 14553 2975 14611 2981
rect 14553 2941 14565 2975
rect 14599 2941 14611 2975
rect 14553 2935 14611 2941
rect 14829 2975 14887 2981
rect 14829 2941 14841 2975
rect 14875 2972 14887 2975
rect 15580 2972 15608 3000
rect 14875 2944 15608 2972
rect 14875 2941 14887 2944
rect 14829 2935 14887 2941
rect 14568 2904 14596 2935
rect 14642 2904 14648 2916
rect 14568 2876 14648 2904
rect 14642 2864 14648 2876
rect 14700 2864 14706 2916
rect 12768 2808 13308 2836
rect 12768 2796 12774 2808
rect 13814 2796 13820 2848
rect 13872 2836 13878 2848
rect 13909 2839 13967 2845
rect 13909 2836 13921 2839
rect 13872 2808 13921 2836
rect 13872 2796 13878 2808
rect 13909 2805 13921 2808
rect 13955 2836 13967 2839
rect 14182 2836 14188 2848
rect 13955 2808 14188 2836
rect 13955 2805 13967 2808
rect 13909 2799 13967 2805
rect 14182 2796 14188 2808
rect 14240 2796 14246 2848
rect 552 2746 15520 2768
rect 552 2694 4100 2746
rect 4152 2694 4164 2746
rect 4216 2694 4228 2746
rect 4280 2694 4292 2746
rect 4344 2694 4356 2746
rect 4408 2694 7802 2746
rect 7854 2694 7866 2746
rect 7918 2694 7930 2746
rect 7982 2694 7994 2746
rect 8046 2694 8058 2746
rect 8110 2694 11504 2746
rect 11556 2694 11568 2746
rect 11620 2694 11632 2746
rect 11684 2694 11696 2746
rect 11748 2694 11760 2746
rect 11812 2694 15206 2746
rect 15258 2694 15270 2746
rect 15322 2694 15334 2746
rect 15386 2694 15398 2746
rect 15450 2694 15462 2746
rect 15514 2694 15520 2746
rect 552 2672 15520 2694
rect 2317 2635 2375 2641
rect 2317 2601 2329 2635
rect 2363 2632 2375 2635
rect 3050 2632 3056 2644
rect 2363 2604 3056 2632
rect 2363 2601 2375 2604
rect 2317 2595 2375 2601
rect 3050 2592 3056 2604
rect 3108 2592 3114 2644
rect 3142 2592 3148 2644
rect 3200 2632 3206 2644
rect 3200 2604 4752 2632
rect 3200 2592 3206 2604
rect 3142 2505 3148 2508
rect 3120 2499 3148 2505
rect 3120 2465 3132 2499
rect 3120 2459 3148 2465
rect 3142 2456 3148 2459
rect 3200 2456 3206 2508
rect 3234 2456 3240 2508
rect 3292 2456 3298 2508
rect 4019 2499 4077 2505
rect 4019 2496 4031 2499
rect 3896 2468 4031 2496
rect 3896 2440 3924 2468
rect 4019 2465 4031 2468
rect 4065 2465 4077 2499
rect 4724 2496 4752 2604
rect 5902 2592 5908 2644
rect 5960 2632 5966 2644
rect 6457 2635 6515 2641
rect 6457 2632 6469 2635
rect 5960 2604 6469 2632
rect 5960 2592 5966 2604
rect 6457 2601 6469 2604
rect 6503 2601 6515 2635
rect 6457 2595 6515 2601
rect 6656 2604 8156 2632
rect 6546 2524 6552 2576
rect 6604 2524 6610 2576
rect 6656 2496 6684 2604
rect 7561 2567 7619 2573
rect 7561 2533 7573 2567
rect 7607 2564 7619 2567
rect 7742 2564 7748 2576
rect 7607 2536 7748 2564
rect 7607 2533 7619 2536
rect 7561 2527 7619 2533
rect 7742 2524 7748 2536
rect 7800 2524 7806 2576
rect 4724 2468 6684 2496
rect 4019 2459 4077 2465
rect 7282 2456 7288 2508
rect 7340 2496 7346 2508
rect 8128 2505 8156 2604
rect 10870 2592 10876 2644
rect 10928 2632 10934 2644
rect 11609 2635 11667 2641
rect 11609 2632 11621 2635
rect 10928 2604 11621 2632
rect 10928 2592 10934 2604
rect 11609 2601 11621 2604
rect 11655 2632 11667 2635
rect 12710 2632 12716 2644
rect 11655 2604 12716 2632
rect 11655 2601 11667 2604
rect 11609 2595 11667 2601
rect 12710 2592 12716 2604
rect 12768 2592 12774 2644
rect 12986 2592 12992 2644
rect 13044 2592 13050 2644
rect 13173 2635 13231 2641
rect 13173 2601 13185 2635
rect 13219 2632 13231 2635
rect 14090 2632 14096 2644
rect 13219 2604 14096 2632
rect 13219 2601 13231 2604
rect 13173 2595 13231 2601
rect 14090 2592 14096 2604
rect 14148 2592 14154 2644
rect 8294 2524 8300 2576
rect 8352 2524 8358 2576
rect 13004 2564 13032 2592
rect 14550 2564 14556 2576
rect 10612 2536 11376 2564
rect 13004 2536 14556 2564
rect 10612 2508 10640 2536
rect 7377 2499 7435 2505
rect 7377 2496 7389 2499
rect 7340 2468 7389 2496
rect 7340 2456 7346 2468
rect 7377 2465 7389 2468
rect 7423 2465 7435 2499
rect 7377 2459 7435 2465
rect 8113 2499 8171 2505
rect 8113 2465 8125 2499
rect 8159 2496 8171 2499
rect 8478 2496 8484 2508
rect 8159 2468 8484 2496
rect 8159 2465 8171 2468
rect 8113 2459 8171 2465
rect 8478 2456 8484 2468
rect 8536 2456 8542 2508
rect 10594 2456 10600 2508
rect 10652 2456 10658 2508
rect 10686 2456 10692 2508
rect 10744 2456 10750 2508
rect 10962 2456 10968 2508
rect 11020 2456 11026 2508
rect 11348 2505 11376 2536
rect 14550 2524 14556 2536
rect 14608 2524 14614 2576
rect 11149 2499 11207 2505
rect 11149 2465 11161 2499
rect 11195 2465 11207 2499
rect 11149 2459 11207 2465
rect 11333 2499 11391 2505
rect 11333 2465 11345 2499
rect 11379 2465 11391 2499
rect 11333 2459 11391 2465
rect 2958 2388 2964 2440
rect 3016 2388 3022 2440
rect 3878 2388 3884 2440
rect 3936 2388 3942 2440
rect 4154 2388 4160 2440
rect 4212 2388 4218 2440
rect 7745 2431 7803 2437
rect 7745 2397 7757 2431
rect 7791 2428 7803 2431
rect 10980 2428 11008 2456
rect 7791 2400 11008 2428
rect 11057 2431 11115 2437
rect 7791 2397 7803 2400
rect 7745 2391 7803 2397
rect 11057 2397 11069 2431
rect 11103 2397 11115 2431
rect 11057 2391 11115 2397
rect 3513 2363 3571 2369
rect 3513 2329 3525 2363
rect 3559 2360 3571 2363
rect 3694 2360 3700 2372
rect 3559 2332 3700 2360
rect 3559 2329 3571 2332
rect 3513 2323 3571 2329
rect 3694 2320 3700 2332
rect 3752 2320 3758 2372
rect 7193 2363 7251 2369
rect 7193 2360 7205 2363
rect 4448 2332 7205 2360
rect 4154 2252 4160 2304
rect 4212 2292 4218 2304
rect 4448 2292 4476 2332
rect 7193 2329 7205 2332
rect 7239 2360 7251 2363
rect 10505 2363 10563 2369
rect 10505 2360 10517 2363
rect 7239 2332 10517 2360
rect 7239 2329 7251 2332
rect 7193 2323 7251 2329
rect 10505 2329 10517 2332
rect 10551 2360 10563 2363
rect 11072 2360 11100 2391
rect 10551 2332 11100 2360
rect 10551 2329 10563 2332
rect 10505 2323 10563 2329
rect 4212 2264 4476 2292
rect 4212 2252 4218 2264
rect 6730 2252 6736 2304
rect 6788 2292 6794 2304
rect 11164 2292 11192 2459
rect 11422 2456 11428 2508
rect 11480 2496 11486 2508
rect 12526 2496 12532 2508
rect 11480 2468 12532 2496
rect 11480 2456 11486 2468
rect 12526 2456 12532 2468
rect 12584 2456 12590 2508
rect 12986 2456 12992 2508
rect 13044 2496 13050 2508
rect 13044 2468 13216 2496
rect 13044 2456 13050 2468
rect 13078 2388 13084 2440
rect 13136 2388 13142 2440
rect 13188 2428 13216 2468
rect 13262 2456 13268 2508
rect 13320 2496 13326 2508
rect 13633 2499 13691 2505
rect 13633 2496 13645 2499
rect 13320 2468 13645 2496
rect 13320 2456 13326 2468
rect 13633 2465 13645 2468
rect 13679 2465 13691 2499
rect 14366 2496 14372 2508
rect 13633 2459 13691 2465
rect 13740 2468 14372 2496
rect 13740 2428 13768 2468
rect 14366 2456 14372 2468
rect 14424 2496 14430 2508
rect 14645 2499 14703 2505
rect 14645 2496 14657 2499
rect 14424 2468 14657 2496
rect 14424 2456 14430 2468
rect 14645 2465 14657 2468
rect 14691 2465 14703 2499
rect 14645 2459 14703 2465
rect 13188 2400 13768 2428
rect 13814 2388 13820 2440
rect 13872 2388 13878 2440
rect 14737 2431 14795 2437
rect 14737 2397 14749 2431
rect 14783 2397 14795 2431
rect 14737 2391 14795 2397
rect 12894 2320 12900 2372
rect 12952 2320 12958 2372
rect 13096 2360 13124 2388
rect 14458 2360 14464 2372
rect 13096 2332 14464 2360
rect 14458 2320 14464 2332
rect 14516 2360 14522 2372
rect 14752 2360 14780 2391
rect 14516 2332 14780 2360
rect 14516 2320 14522 2332
rect 11514 2292 11520 2304
rect 6788 2264 11520 2292
rect 6788 2252 6794 2264
rect 11514 2252 11520 2264
rect 11572 2252 11578 2304
rect 12912 2292 12940 2320
rect 13541 2295 13599 2301
rect 13541 2292 13553 2295
rect 12912 2264 13553 2292
rect 13541 2261 13553 2264
rect 13587 2261 13599 2295
rect 13541 2255 13599 2261
rect 14182 2252 14188 2304
rect 14240 2252 14246 2304
rect 552 2202 15364 2224
rect 552 2150 2249 2202
rect 2301 2150 2313 2202
rect 2365 2150 2377 2202
rect 2429 2150 2441 2202
rect 2493 2150 2505 2202
rect 2557 2150 5951 2202
rect 6003 2150 6015 2202
rect 6067 2150 6079 2202
rect 6131 2150 6143 2202
rect 6195 2150 6207 2202
rect 6259 2150 9653 2202
rect 9705 2150 9717 2202
rect 9769 2150 9781 2202
rect 9833 2150 9845 2202
rect 9897 2150 9909 2202
rect 9961 2150 13355 2202
rect 13407 2150 13419 2202
rect 13471 2150 13483 2202
rect 13535 2150 13547 2202
rect 13599 2150 13611 2202
rect 13663 2150 15364 2202
rect 552 2128 15364 2150
rect 4433 2091 4491 2097
rect 4433 2057 4445 2091
rect 4479 2088 4491 2091
rect 4890 2088 4896 2100
rect 4479 2060 4896 2088
rect 4479 2057 4491 2060
rect 4433 2051 4491 2057
rect 4890 2048 4896 2060
rect 4948 2048 4954 2100
rect 8662 2088 8668 2100
rect 5552 2060 8668 2088
rect 3234 1912 3240 1964
rect 3292 1952 3298 1964
rect 3513 1955 3571 1961
rect 3513 1952 3525 1955
rect 3292 1924 3525 1952
rect 3292 1912 3298 1924
rect 3513 1921 3525 1924
rect 3559 1921 3571 1955
rect 5077 1955 5135 1961
rect 5077 1952 5089 1955
rect 3513 1915 3571 1921
rect 4356 1924 5089 1952
rect 3605 1887 3663 1893
rect 3605 1853 3617 1887
rect 3651 1884 3663 1887
rect 4154 1884 4160 1896
rect 3651 1856 4160 1884
rect 3651 1853 3663 1856
rect 3605 1847 3663 1853
rect 4154 1844 4160 1856
rect 4212 1844 4218 1896
rect 2958 1776 2964 1828
rect 3016 1816 3022 1828
rect 4356 1816 4384 1924
rect 5077 1921 5089 1924
rect 5123 1952 5135 1955
rect 5552 1952 5580 2060
rect 8662 2048 8668 2060
rect 8720 2048 8726 2100
rect 9033 2091 9091 2097
rect 9033 2057 9045 2091
rect 9079 2088 9091 2091
rect 9490 2088 9496 2100
rect 9079 2060 9496 2088
rect 9079 2057 9091 2060
rect 9033 2051 9091 2057
rect 9490 2048 9496 2060
rect 9548 2048 9554 2100
rect 10686 2048 10692 2100
rect 10744 2088 10750 2100
rect 10965 2091 11023 2097
rect 10965 2088 10977 2091
rect 10744 2060 10977 2088
rect 10744 2048 10750 2060
rect 10965 2057 10977 2060
rect 11011 2057 11023 2091
rect 10965 2051 11023 2057
rect 11514 2048 11520 2100
rect 11572 2088 11578 2100
rect 12802 2088 12808 2100
rect 11572 2060 12808 2088
rect 11572 2048 11578 2060
rect 12802 2048 12808 2060
rect 12860 2048 12866 2100
rect 13170 2048 13176 2100
rect 13228 2048 13234 2100
rect 14645 2091 14703 2097
rect 14645 2057 14657 2091
rect 14691 2088 14703 2091
rect 15562 2088 15568 2100
rect 14691 2060 15568 2088
rect 14691 2057 14703 2060
rect 14645 2051 14703 2057
rect 15562 2048 15568 2060
rect 15620 2048 15626 2100
rect 5626 1980 5632 2032
rect 5684 1980 5690 2032
rect 6362 2020 6368 2032
rect 5828 1992 6368 2020
rect 5123 1924 5580 1952
rect 5644 1952 5672 1980
rect 5828 1952 5856 1992
rect 6362 1980 6368 1992
rect 6420 1980 6426 2032
rect 7190 1980 7196 2032
rect 7248 2020 7254 2032
rect 8754 2020 8760 2032
rect 7248 1992 8760 2020
rect 7248 1980 7254 1992
rect 8754 1980 8760 1992
rect 8812 2020 8818 2032
rect 13078 2020 13084 2032
rect 8812 1992 9812 2020
rect 8812 1980 8818 1992
rect 5644 1924 5856 1952
rect 5123 1921 5135 1924
rect 5077 1915 5135 1921
rect 6086 1912 6092 1964
rect 6144 1952 6150 1964
rect 6822 1952 6828 1964
rect 6144 1924 6828 1952
rect 6144 1912 6150 1924
rect 6822 1912 6828 1924
rect 6880 1912 6886 1964
rect 8036 1924 8616 1952
rect 5258 1893 5264 1896
rect 5236 1887 5264 1893
rect 5236 1853 5248 1887
rect 5236 1847 5264 1853
rect 5258 1844 5264 1847
rect 5316 1844 5322 1896
rect 5350 1844 5356 1896
rect 5408 1844 5414 1896
rect 6178 1844 6184 1896
rect 6236 1884 6242 1896
rect 6273 1887 6331 1893
rect 6273 1884 6285 1887
rect 6236 1856 6285 1884
rect 6236 1844 6242 1856
rect 6273 1853 6285 1856
rect 6319 1884 6331 1887
rect 6730 1884 6736 1896
rect 6319 1856 6736 1884
rect 6319 1853 6331 1856
rect 6273 1847 6331 1853
rect 6730 1844 6736 1856
rect 6788 1844 6794 1896
rect 3016 1788 4384 1816
rect 3016 1776 3022 1788
rect 3234 1708 3240 1760
rect 3292 1708 3298 1760
rect 5258 1708 5264 1760
rect 5316 1748 5322 1760
rect 7742 1748 7748 1760
rect 5316 1720 7748 1748
rect 5316 1708 5322 1720
rect 7742 1708 7748 1720
rect 7800 1748 7806 1760
rect 8036 1757 8064 1924
rect 8478 1844 8484 1896
rect 8536 1844 8542 1896
rect 8588 1893 8616 1924
rect 8573 1887 8631 1893
rect 8573 1853 8585 1887
rect 8619 1853 8631 1887
rect 8573 1847 8631 1853
rect 8662 1844 8668 1896
rect 8720 1884 8726 1896
rect 8757 1887 8815 1893
rect 8757 1884 8769 1887
rect 8720 1856 8769 1884
rect 8720 1844 8726 1856
rect 8757 1853 8769 1856
rect 8803 1884 8815 1887
rect 9214 1884 9220 1896
rect 8803 1856 9220 1884
rect 8803 1853 8815 1856
rect 8757 1847 8815 1853
rect 9214 1844 9220 1856
rect 9272 1844 9278 1896
rect 9784 1893 9812 1992
rect 12360 1992 13084 2020
rect 9953 1955 10011 1961
rect 9953 1921 9965 1955
rect 9999 1952 10011 1955
rect 10134 1952 10140 1964
rect 9999 1924 10140 1952
rect 9999 1921 10011 1924
rect 9953 1915 10011 1921
rect 10134 1912 10140 1924
rect 10192 1912 10198 1964
rect 10226 1912 10232 1964
rect 10284 1912 10290 1964
rect 11146 1912 11152 1964
rect 11204 1952 11210 1964
rect 12360 1961 12388 1992
rect 13078 1980 13084 1992
rect 13136 1980 13142 2032
rect 11517 1955 11575 1961
rect 11517 1952 11529 1955
rect 11204 1924 11529 1952
rect 11204 1912 11210 1924
rect 11517 1921 11529 1924
rect 11563 1952 11575 1955
rect 12345 1955 12403 1961
rect 12345 1952 12357 1955
rect 11563 1924 12357 1952
rect 11563 1921 11575 1924
rect 11517 1915 11575 1921
rect 12345 1921 12357 1924
rect 12391 1921 12403 1955
rect 12345 1915 12403 1921
rect 12434 1912 12440 1964
rect 12492 1912 12498 1964
rect 13188 1952 13216 2048
rect 13354 1980 13360 2032
rect 13412 2020 13418 2032
rect 13630 2020 13636 2032
rect 13412 1992 13636 2020
rect 13412 1980 13418 1992
rect 13630 1980 13636 1992
rect 13688 2020 13694 2032
rect 14093 2023 14151 2029
rect 14093 2020 14105 2023
rect 13688 1992 14105 2020
rect 13688 1980 13694 1992
rect 14093 1989 14105 1992
rect 14139 1989 14151 2023
rect 14093 1983 14151 1989
rect 15010 1980 15016 2032
rect 15068 1980 15074 2032
rect 13188 1924 14596 1952
rect 9769 1887 9827 1893
rect 9769 1853 9781 1887
rect 9815 1853 9827 1887
rect 9769 1847 9827 1853
rect 9861 1887 9919 1893
rect 9861 1853 9873 1887
rect 9907 1884 9919 1887
rect 10244 1884 10272 1912
rect 9907 1856 10272 1884
rect 9907 1853 9919 1856
rect 9861 1847 9919 1853
rect 11238 1844 11244 1896
rect 11296 1844 11302 1896
rect 11425 1887 11483 1893
rect 11425 1853 11437 1887
rect 11471 1884 11483 1887
rect 12452 1884 12480 1912
rect 11471 1856 12480 1884
rect 11471 1853 11483 1856
rect 11425 1847 11483 1853
rect 14182 1844 14188 1896
rect 14240 1884 14246 1896
rect 14568 1893 14596 1924
rect 14277 1887 14335 1893
rect 14277 1884 14289 1887
rect 14240 1856 14289 1884
rect 14240 1844 14246 1856
rect 14277 1853 14289 1856
rect 14323 1853 14335 1887
rect 14277 1847 14335 1853
rect 14553 1887 14611 1893
rect 14553 1853 14565 1887
rect 14599 1853 14611 1887
rect 14553 1847 14611 1853
rect 14829 1887 14887 1893
rect 14829 1853 14841 1887
rect 14875 1884 14887 1887
rect 15028 1884 15056 1980
rect 14875 1856 15056 1884
rect 14875 1853 14887 1856
rect 14829 1847 14887 1853
rect 8113 1819 8171 1825
rect 8113 1785 8125 1819
rect 8159 1816 8171 1819
rect 8159 1788 9444 1816
rect 8159 1785 8171 1788
rect 8113 1779 8171 1785
rect 9416 1757 9444 1788
rect 10042 1776 10048 1828
rect 10100 1776 10106 1828
rect 11256 1816 11284 1844
rect 12161 1819 12219 1825
rect 12161 1816 12173 1819
rect 11256 1788 12173 1816
rect 12161 1785 12173 1788
rect 12207 1816 12219 1819
rect 12434 1816 12440 1828
rect 12207 1788 12440 1816
rect 12207 1785 12219 1788
rect 12161 1779 12219 1785
rect 12434 1776 12440 1788
rect 12492 1776 12498 1828
rect 12710 1776 12716 1828
rect 12768 1776 12774 1828
rect 12986 1776 12992 1828
rect 13044 1816 13050 1828
rect 13044 1788 14412 1816
rect 13044 1776 13050 1788
rect 8021 1751 8079 1757
rect 8021 1748 8033 1751
rect 7800 1720 8033 1748
rect 7800 1708 7806 1720
rect 8021 1717 8033 1720
rect 8067 1717 8079 1751
rect 8021 1711 8079 1717
rect 9401 1751 9459 1757
rect 9401 1717 9413 1751
rect 9447 1717 9459 1751
rect 10060 1748 10088 1776
rect 11333 1751 11391 1757
rect 11333 1748 11345 1751
rect 10060 1720 11345 1748
rect 9401 1711 9459 1717
rect 11333 1717 11345 1720
rect 11379 1748 11391 1751
rect 11422 1748 11428 1760
rect 11379 1720 11428 1748
rect 11379 1717 11391 1720
rect 11333 1711 11391 1717
rect 11422 1708 11428 1720
rect 11480 1708 11486 1760
rect 11793 1751 11851 1757
rect 11793 1717 11805 1751
rect 11839 1748 11851 1751
rect 11882 1748 11888 1760
rect 11839 1720 11888 1748
rect 11839 1717 11851 1720
rect 11793 1711 11851 1717
rect 11882 1708 11888 1720
rect 11940 1708 11946 1760
rect 12066 1708 12072 1760
rect 12124 1748 12130 1760
rect 12253 1751 12311 1757
rect 12253 1748 12265 1751
rect 12124 1720 12265 1748
rect 12124 1708 12130 1720
rect 12253 1717 12265 1720
rect 12299 1748 12311 1751
rect 13998 1748 14004 1760
rect 12299 1720 14004 1748
rect 12299 1717 12311 1720
rect 12253 1711 12311 1717
rect 13998 1708 14004 1720
rect 14056 1708 14062 1760
rect 14384 1757 14412 1788
rect 14369 1751 14427 1757
rect 14369 1717 14381 1751
rect 14415 1717 14427 1751
rect 14369 1711 14427 1717
rect 552 1658 15520 1680
rect 552 1606 4100 1658
rect 4152 1606 4164 1658
rect 4216 1606 4228 1658
rect 4280 1606 4292 1658
rect 4344 1606 4356 1658
rect 4408 1606 7802 1658
rect 7854 1606 7866 1658
rect 7918 1606 7930 1658
rect 7982 1606 7994 1658
rect 8046 1606 8058 1658
rect 8110 1606 11504 1658
rect 11556 1606 11568 1658
rect 11620 1606 11632 1658
rect 11684 1606 11696 1658
rect 11748 1606 11760 1658
rect 11812 1606 15206 1658
rect 15258 1606 15270 1658
rect 15322 1606 15334 1658
rect 15386 1606 15398 1658
rect 15450 1606 15462 1658
rect 15514 1606 15520 1658
rect 552 1584 15520 1606
rect 3142 1504 3148 1556
rect 3200 1504 3206 1556
rect 3786 1504 3792 1556
rect 3844 1504 3850 1556
rect 5258 1544 5264 1556
rect 4632 1516 5264 1544
rect 3160 1476 3188 1504
rect 2884 1448 3188 1476
rect 2774 1368 2780 1420
rect 2832 1368 2838 1420
rect 2884 1349 2912 1448
rect 4632 1417 4660 1516
rect 5258 1504 5264 1516
rect 5316 1504 5322 1556
rect 6181 1547 6239 1553
rect 6181 1513 6193 1547
rect 6227 1544 6239 1547
rect 6270 1544 6276 1556
rect 6227 1516 6276 1544
rect 6227 1513 6239 1516
rect 6181 1507 6239 1513
rect 6270 1504 6276 1516
rect 6328 1504 6334 1556
rect 6914 1504 6920 1556
rect 6972 1544 6978 1556
rect 7009 1547 7067 1553
rect 7009 1544 7021 1547
rect 6972 1516 7021 1544
rect 6972 1504 6978 1516
rect 7009 1513 7021 1516
rect 7055 1513 7067 1547
rect 7009 1507 7067 1513
rect 7377 1547 7435 1553
rect 7377 1513 7389 1547
rect 7423 1544 7435 1547
rect 7466 1544 7472 1556
rect 7423 1516 7472 1544
rect 7423 1513 7435 1516
rect 7377 1507 7435 1513
rect 7466 1504 7472 1516
rect 7524 1504 7530 1556
rect 11882 1504 11888 1556
rect 11940 1504 11946 1556
rect 12529 1547 12587 1553
rect 12529 1513 12541 1547
rect 12575 1544 12587 1547
rect 12710 1544 12716 1556
rect 12575 1516 12716 1544
rect 12575 1513 12587 1516
rect 12529 1507 12587 1513
rect 12710 1504 12716 1516
rect 12768 1504 12774 1556
rect 12802 1504 12808 1556
rect 12860 1544 12866 1556
rect 12860 1516 13124 1544
rect 12860 1504 12866 1516
rect 5350 1476 5356 1488
rect 4724 1448 5356 1476
rect 3421 1411 3479 1417
rect 3421 1408 3433 1411
rect 3160 1380 3433 1408
rect 3160 1349 3188 1380
rect 3421 1377 3433 1380
rect 3467 1377 3479 1411
rect 3421 1371 3479 1377
rect 4617 1411 4675 1417
rect 4617 1377 4629 1411
rect 4663 1377 4675 1411
rect 4617 1371 4675 1377
rect 2869 1343 2927 1349
rect 2869 1309 2881 1343
rect 2915 1309 2927 1343
rect 2869 1303 2927 1309
rect 3145 1343 3203 1349
rect 3145 1309 3157 1343
rect 3191 1309 3203 1343
rect 3145 1303 3203 1309
rect 3234 1300 3240 1352
rect 3292 1340 3298 1352
rect 4724 1349 4752 1448
rect 5350 1436 5356 1448
rect 5408 1436 5414 1488
rect 7558 1436 7564 1488
rect 7616 1476 7622 1488
rect 11517 1479 11575 1485
rect 7616 1448 8156 1476
rect 7616 1436 7622 1448
rect 5261 1411 5319 1417
rect 5261 1377 5273 1411
rect 5307 1408 5319 1411
rect 6086 1408 6092 1420
rect 5307 1380 6092 1408
rect 5307 1377 5319 1380
rect 5261 1371 5319 1377
rect 6086 1368 6092 1380
rect 6144 1368 6150 1420
rect 6549 1411 6607 1417
rect 6549 1377 6561 1411
rect 6595 1408 6607 1411
rect 7190 1408 7196 1420
rect 6595 1380 7196 1408
rect 6595 1377 6607 1380
rect 6549 1371 6607 1377
rect 7190 1368 7196 1380
rect 7248 1368 7254 1420
rect 3329 1343 3387 1349
rect 3329 1340 3341 1343
rect 3292 1312 3341 1340
rect 3292 1300 3298 1312
rect 3329 1309 3341 1312
rect 3375 1309 3387 1343
rect 3329 1303 3387 1309
rect 4709 1343 4767 1349
rect 4709 1309 4721 1343
rect 4755 1309 4767 1343
rect 4709 1303 4767 1309
rect 5353 1343 5411 1349
rect 5353 1309 5365 1343
rect 5399 1340 5411 1343
rect 6178 1340 6184 1352
rect 5399 1312 6184 1340
rect 5399 1309 5411 1312
rect 5353 1303 5411 1309
rect 6178 1300 6184 1312
rect 6236 1300 6242 1352
rect 6638 1300 6644 1352
rect 6696 1300 6702 1352
rect 6825 1343 6883 1349
rect 6825 1309 6837 1343
rect 6871 1340 6883 1343
rect 7006 1340 7012 1352
rect 6871 1312 7012 1340
rect 6871 1309 6883 1312
rect 6825 1303 6883 1309
rect 7006 1300 7012 1312
rect 7064 1300 7070 1352
rect 7466 1300 7472 1352
rect 7524 1300 7530 1352
rect 8128 1349 8156 1448
rect 11517 1445 11529 1479
rect 11563 1476 11575 1479
rect 11900 1476 11928 1504
rect 11563 1448 11928 1476
rect 11563 1445 11575 1448
rect 11517 1439 11575 1445
rect 12250 1436 12256 1488
rect 12308 1476 12314 1488
rect 12986 1476 12992 1488
rect 12308 1448 12992 1476
rect 12308 1436 12314 1448
rect 12986 1436 12992 1448
rect 13044 1436 13050 1488
rect 13096 1476 13124 1516
rect 13262 1504 13268 1556
rect 13320 1544 13326 1556
rect 13357 1547 13415 1553
rect 13357 1544 13369 1547
rect 13320 1516 13369 1544
rect 13320 1504 13326 1516
rect 13357 1513 13369 1516
rect 13403 1513 13415 1547
rect 13357 1507 13415 1513
rect 13722 1504 13728 1556
rect 13780 1504 13786 1556
rect 14366 1504 14372 1556
rect 14424 1504 14430 1556
rect 14642 1504 14648 1556
rect 14700 1504 14706 1556
rect 14734 1504 14740 1556
rect 14792 1504 14798 1556
rect 13541 1479 13599 1485
rect 13541 1476 13553 1479
rect 13096 1448 13553 1476
rect 13541 1445 13553 1448
rect 13587 1445 13599 1479
rect 13541 1439 13599 1445
rect 8205 1411 8263 1417
rect 8205 1377 8217 1411
rect 8251 1408 8263 1411
rect 8662 1408 8668 1420
rect 8251 1380 8668 1408
rect 8251 1377 8263 1380
rect 8205 1371 8263 1377
rect 8662 1368 8668 1380
rect 8720 1368 8726 1420
rect 10502 1368 10508 1420
rect 10560 1368 10566 1420
rect 12897 1411 12955 1417
rect 12897 1408 12909 1411
rect 12176 1380 12909 1408
rect 7561 1343 7619 1349
rect 7561 1309 7573 1343
rect 7607 1309 7619 1343
rect 7561 1303 7619 1309
rect 8113 1343 8171 1349
rect 8113 1309 8125 1343
rect 8159 1309 8171 1343
rect 8113 1303 8171 1309
rect 4985 1275 5043 1281
rect 4985 1241 4997 1275
rect 5031 1272 5043 1275
rect 5718 1272 5724 1284
rect 5031 1244 5724 1272
rect 5031 1241 5043 1244
rect 4985 1235 5043 1241
rect 5718 1232 5724 1244
rect 5776 1232 5782 1284
rect 7024 1272 7052 1300
rect 7576 1272 7604 1303
rect 10594 1300 10600 1352
rect 10652 1300 10658 1352
rect 11422 1300 11428 1352
rect 11480 1340 11486 1352
rect 12176 1340 12204 1380
rect 12897 1377 12909 1380
rect 12943 1377 12955 1411
rect 13740 1408 13768 1504
rect 14553 1411 14611 1417
rect 13740 1380 14504 1408
rect 12897 1371 12955 1377
rect 11480 1312 12204 1340
rect 11480 1300 11486 1312
rect 13078 1300 13084 1352
rect 13136 1300 13142 1352
rect 13170 1300 13176 1352
rect 13228 1340 13234 1352
rect 13725 1343 13783 1349
rect 13725 1340 13737 1343
rect 13228 1312 13737 1340
rect 13228 1300 13234 1312
rect 13725 1309 13737 1312
rect 13771 1309 13783 1343
rect 14476 1340 14504 1380
rect 14553 1377 14565 1411
rect 14599 1408 14611 1411
rect 14752 1408 14780 1504
rect 14599 1380 14780 1408
rect 14829 1411 14887 1417
rect 14599 1377 14611 1380
rect 14553 1371 14611 1377
rect 14829 1377 14841 1411
rect 14875 1377 14887 1411
rect 14829 1371 14887 1377
rect 14844 1340 14872 1371
rect 14476 1312 14872 1340
rect 13725 1303 13783 1309
rect 11333 1275 11391 1281
rect 11333 1272 11345 1275
rect 7024 1244 7604 1272
rect 8404 1244 11345 1272
rect 8404 1216 8432 1244
rect 11333 1241 11345 1244
rect 11379 1272 11391 1275
rect 13906 1272 13912 1284
rect 11379 1244 13912 1272
rect 11379 1241 11391 1244
rect 11333 1235 11391 1241
rect 13906 1232 13912 1244
rect 13964 1232 13970 1284
rect 5626 1164 5632 1216
rect 5684 1164 5690 1216
rect 8386 1164 8392 1216
rect 8444 1164 8450 1216
rect 8478 1164 8484 1216
rect 8536 1164 8542 1216
rect 10134 1164 10140 1216
rect 10192 1164 10198 1216
rect 552 1114 15364 1136
rect 552 1062 2249 1114
rect 2301 1062 2313 1114
rect 2365 1062 2377 1114
rect 2429 1062 2441 1114
rect 2493 1062 2505 1114
rect 2557 1062 5951 1114
rect 6003 1062 6015 1114
rect 6067 1062 6079 1114
rect 6131 1062 6143 1114
rect 6195 1062 6207 1114
rect 6259 1062 9653 1114
rect 9705 1062 9717 1114
rect 9769 1062 9781 1114
rect 9833 1062 9845 1114
rect 9897 1062 9909 1114
rect 9961 1062 13355 1114
rect 13407 1062 13419 1114
rect 13471 1062 13483 1114
rect 13535 1062 13547 1114
rect 13599 1062 13611 1114
rect 13663 1062 15364 1114
rect 552 1040 15364 1062
rect 1118 960 1124 1012
rect 1176 960 1182 1012
rect 3418 960 3424 1012
rect 3476 960 3482 1012
rect 4157 1003 4215 1009
rect 4157 969 4169 1003
rect 4203 1000 4215 1003
rect 4522 1000 4528 1012
rect 4203 972 4528 1000
rect 4203 969 4215 972
rect 4157 963 4215 969
rect 4522 960 4528 972
rect 4580 960 4586 1012
rect 5074 960 5080 1012
rect 5132 1000 5138 1012
rect 5169 1003 5227 1009
rect 5169 1000 5181 1003
rect 5132 972 5181 1000
rect 5132 960 5138 972
rect 5169 969 5181 972
rect 5215 969 5227 1003
rect 5169 963 5227 969
rect 5626 960 5632 1012
rect 5684 960 5690 1012
rect 5718 960 5724 1012
rect 5776 960 5782 1012
rect 6273 1003 6331 1009
rect 6273 969 6285 1003
rect 6319 1000 6331 1003
rect 6638 1000 6644 1012
rect 6319 972 6644 1000
rect 6319 969 6331 972
rect 6273 963 6331 969
rect 6638 960 6644 972
rect 6696 960 6702 1012
rect 7190 960 7196 1012
rect 7248 960 7254 1012
rect 7650 960 7656 1012
rect 7708 1000 7714 1012
rect 8021 1003 8079 1009
rect 8021 1000 8033 1003
rect 7708 972 8033 1000
rect 7708 960 7714 972
rect 8021 969 8033 972
rect 8067 969 8079 1003
rect 8021 963 8079 969
rect 8478 960 8484 1012
rect 8536 960 8542 1012
rect 9677 1003 9735 1009
rect 9677 969 9689 1003
rect 9723 1000 9735 1003
rect 10042 1000 10048 1012
rect 9723 972 10048 1000
rect 9723 969 9735 972
rect 9677 963 9735 969
rect 10042 960 10048 972
rect 10100 960 10106 1012
rect 10134 960 10140 1012
rect 10192 960 10198 1012
rect 10229 1003 10287 1009
rect 10229 969 10241 1003
rect 10275 1000 10287 1003
rect 10318 1000 10324 1012
rect 10275 972 10324 1000
rect 10275 969 10287 972
rect 10229 963 10287 969
rect 10318 960 10324 972
rect 10376 960 10382 1012
rect 11241 1003 11299 1009
rect 11241 969 11253 1003
rect 11287 1000 11299 1003
rect 11330 1000 11336 1012
rect 11287 972 11336 1000
rect 11287 969 11299 972
rect 11241 963 11299 969
rect 11330 960 11336 972
rect 11388 960 11394 1012
rect 12253 1003 12311 1009
rect 12253 969 12265 1003
rect 12299 1000 12311 1003
rect 12342 1000 12348 1012
rect 12299 972 12348 1000
rect 12299 969 12311 972
rect 12253 963 12311 969
rect 12342 960 12348 972
rect 12400 960 12406 1012
rect 12434 960 12440 1012
rect 12492 1000 12498 1012
rect 13265 1003 13323 1009
rect 13265 1000 13277 1003
rect 12492 972 13277 1000
rect 12492 960 12498 972
rect 13265 969 13277 972
rect 13311 969 13323 1003
rect 13265 963 13323 969
rect 13814 960 13820 1012
rect 13872 1000 13878 1012
rect 14185 1003 14243 1009
rect 14185 1000 14197 1003
rect 13872 972 14197 1000
rect 13872 960 13878 972
rect 14185 969 14197 972
rect 14231 969 14243 1003
rect 14185 963 14243 969
rect 14550 960 14556 1012
rect 14608 1000 14614 1012
rect 14829 1003 14887 1009
rect 14829 1000 14841 1003
rect 14608 972 14841 1000
rect 14608 960 14614 972
rect 14829 969 14841 972
rect 14875 969 14887 1003
rect 14829 963 14887 969
rect 2133 935 2191 941
rect 2133 901 2145 935
rect 2179 932 2191 935
rect 4706 932 4712 944
rect 2179 904 4712 932
rect 2179 901 2191 904
rect 2133 895 2191 901
rect 4706 892 4712 904
rect 4764 892 4770 944
rect 2774 824 2780 876
rect 2832 824 2838 876
rect 934 756 940 808
rect 992 756 998 808
rect 1946 756 1952 808
rect 2004 756 2010 808
rect 2792 728 2820 824
rect 2866 756 2872 808
rect 2924 796 2930 808
rect 3237 799 3295 805
rect 3237 796 3249 799
rect 2924 768 3249 796
rect 2924 756 2930 768
rect 3237 765 3249 768
rect 3283 765 3295 799
rect 3237 759 3295 765
rect 3970 756 3976 808
rect 4028 756 4034 808
rect 4982 756 4988 808
rect 5040 756 5046 808
rect 5644 796 5672 960
rect 5736 864 5764 960
rect 5905 867 5963 873
rect 5905 864 5917 867
rect 5736 836 5917 864
rect 5905 833 5917 836
rect 5951 833 5963 867
rect 8386 864 8392 876
rect 5905 827 5963 833
rect 6564 836 8392 864
rect 5997 799 6055 805
rect 5997 796 6009 799
rect 5644 768 6009 796
rect 5997 765 6009 768
rect 6043 765 6055 799
rect 5997 759 6055 765
rect 6178 756 6184 808
rect 6236 796 6242 808
rect 6457 799 6515 805
rect 6457 796 6469 799
rect 6236 768 6469 796
rect 6236 756 6242 768
rect 6457 765 6469 768
rect 6503 765 6515 799
rect 6457 759 6515 765
rect 6564 728 6592 836
rect 8386 824 8392 836
rect 8444 824 8450 876
rect 8496 864 8524 960
rect 9125 867 9183 873
rect 9125 864 9137 867
rect 8496 836 9137 864
rect 9125 833 9137 836
rect 9171 833 9183 867
rect 10152 864 10180 960
rect 13906 892 13912 944
rect 13964 892 13970 944
rect 9125 827 9183 833
rect 9232 836 10180 864
rect 13924 864 13952 892
rect 14093 867 14151 873
rect 14093 864 14105 867
rect 13924 836 14105 864
rect 7006 756 7012 808
rect 7064 756 7070 808
rect 7374 756 7380 808
rect 7432 756 7438 808
rect 7466 756 7472 808
rect 7524 756 7530 808
rect 8202 756 8208 808
rect 8260 756 8266 808
rect 9232 805 9260 836
rect 14093 833 14105 836
rect 14139 833 14151 867
rect 14093 827 14151 833
rect 9217 799 9275 805
rect 9217 765 9229 799
rect 9263 765 9275 799
rect 9217 759 9275 765
rect 9493 799 9551 805
rect 9493 765 9505 799
rect 9539 765 9551 799
rect 9493 759 9551 765
rect 7392 728 7420 756
rect 2792 700 6592 728
rect 6656 700 7420 728
rect 6656 669 6684 700
rect 6641 663 6699 669
rect 6641 629 6653 663
rect 6687 629 6699 663
rect 7484 660 7512 756
rect 8938 688 8944 740
rect 8996 728 9002 740
rect 9508 728 9536 759
rect 10042 756 10048 808
rect 10100 756 10106 808
rect 10502 756 10508 808
rect 10560 756 10566 808
rect 11054 756 11060 808
rect 11112 756 11118 808
rect 12066 756 12072 808
rect 12124 756 12130 808
rect 13078 756 13084 808
rect 13136 756 13142 808
rect 13722 756 13728 808
rect 13780 756 13786 808
rect 13909 799 13967 805
rect 13909 765 13921 799
rect 13955 765 13967 799
rect 13909 759 13967 765
rect 8996 700 9536 728
rect 10520 728 10548 756
rect 13924 728 13952 759
rect 13998 756 14004 808
rect 14056 796 14062 808
rect 14369 799 14427 805
rect 14369 796 14381 799
rect 14056 768 14381 796
rect 14056 756 14062 768
rect 14369 765 14381 768
rect 14415 765 14427 799
rect 14369 759 14427 765
rect 15010 756 15016 808
rect 15068 756 15074 808
rect 14918 728 14924 740
rect 10520 700 14924 728
rect 8996 688 9002 700
rect 14918 688 14924 700
rect 14976 688 14982 740
rect 8849 663 8907 669
rect 8849 660 8861 663
rect 7484 632 8861 660
rect 6641 623 6699 629
rect 8849 629 8861 632
rect 8895 629 8907 663
rect 8849 623 8907 629
rect 14553 663 14611 669
rect 14553 629 14565 663
rect 14599 660 14611 663
rect 15102 660 15108 672
rect 14599 632 15108 660
rect 14599 629 14611 632
rect 14553 623 14611 629
rect 15102 620 15108 632
rect 15160 620 15166 672
rect 552 570 15520 592
rect 552 518 4100 570
rect 4152 518 4164 570
rect 4216 518 4228 570
rect 4280 518 4292 570
rect 4344 518 4356 570
rect 4408 518 7802 570
rect 7854 518 7866 570
rect 7918 518 7930 570
rect 7982 518 7994 570
rect 8046 518 8058 570
rect 8110 518 11504 570
rect 11556 518 11568 570
rect 11620 518 11632 570
rect 11684 518 11696 570
rect 11748 518 11760 570
rect 11812 518 15206 570
rect 15258 518 15270 570
rect 15322 518 15334 570
rect 15386 518 15398 570
rect 15450 518 15462 570
rect 15514 518 15520 570
rect 552 496 15520 518
rect 8018 416 8024 468
rect 8076 456 8082 468
rect 8202 456 8208 468
rect 8076 428 8208 456
rect 8076 416 8082 428
rect 8202 416 8208 428
rect 8260 416 8266 468
<< via1 >>
rect 7472 6740 7524 6792
rect 10876 6740 10928 6792
rect 12256 6740 12308 6792
rect 15016 6740 15068 6792
rect 7104 6672 7156 6724
rect 15660 6672 15712 6724
rect 8116 6604 8168 6656
rect 11980 6604 12032 6656
rect 12900 6604 12952 6656
rect 15568 6604 15620 6656
rect 2249 6502 2301 6554
rect 2313 6502 2365 6554
rect 2377 6502 2429 6554
rect 2441 6502 2493 6554
rect 2505 6502 2557 6554
rect 5951 6502 6003 6554
rect 6015 6502 6067 6554
rect 6079 6502 6131 6554
rect 6143 6502 6195 6554
rect 6207 6502 6259 6554
rect 9653 6502 9705 6554
rect 9717 6502 9769 6554
rect 9781 6502 9833 6554
rect 9845 6502 9897 6554
rect 9909 6502 9961 6554
rect 13355 6502 13407 6554
rect 13419 6502 13471 6554
rect 13483 6502 13535 6554
rect 13547 6502 13599 6554
rect 13611 6502 13663 6554
rect 1492 6400 1544 6452
rect 2136 6400 2188 6452
rect 2596 6400 2648 6452
rect 2964 6400 3016 6452
rect 3332 6443 3384 6452
rect 3332 6409 3341 6443
rect 3341 6409 3375 6443
rect 3375 6409 3384 6443
rect 3332 6400 3384 6409
rect 4068 6400 4120 6452
rect 4436 6400 4488 6452
rect 4804 6400 4856 6452
rect 5448 6400 5500 6452
rect 5816 6400 5868 6452
rect 6276 6400 6328 6452
rect 6644 6443 6696 6452
rect 6644 6409 6653 6443
rect 6653 6409 6687 6443
rect 6687 6409 6696 6443
rect 6644 6400 6696 6409
rect 7012 6400 7064 6452
rect 7380 6400 7432 6452
rect 7748 6400 7800 6452
rect 11980 6400 12032 6452
rect 8852 6332 8904 6384
rect 8944 6332 8996 6384
rect 14280 6332 14332 6384
rect 5172 6264 5224 6316
rect 8484 6264 8536 6316
rect 12624 6307 12676 6316
rect 12624 6273 12633 6307
rect 12633 6273 12667 6307
rect 12667 6273 12676 6307
rect 12624 6264 12676 6273
rect 13544 6264 13596 6316
rect 14648 6307 14700 6316
rect 14648 6273 14657 6307
rect 14657 6273 14691 6307
rect 14691 6273 14700 6307
rect 14648 6264 14700 6273
rect 756 6196 808 6248
rect 1308 6196 1360 6248
rect 3608 6196 3660 6248
rect 3884 6196 3936 6248
rect 4528 6196 4580 6248
rect 4712 6239 4764 6248
rect 4712 6205 4721 6239
rect 4721 6205 4755 6239
rect 4755 6205 4764 6239
rect 4712 6196 4764 6205
rect 5356 6239 5408 6248
rect 5356 6205 5365 6239
rect 5365 6205 5399 6239
rect 5399 6205 5408 6239
rect 5356 6196 5408 6205
rect 4988 6128 5040 6180
rect 6184 6239 6236 6248
rect 6184 6205 6193 6239
rect 6193 6205 6227 6239
rect 6227 6205 6236 6239
rect 6184 6196 6236 6205
rect 6828 6239 6880 6248
rect 6828 6205 6837 6239
rect 6837 6205 6871 6239
rect 6871 6205 6880 6239
rect 6828 6196 6880 6205
rect 7380 6239 7432 6248
rect 7380 6205 7389 6239
rect 7389 6205 7423 6239
rect 7423 6205 7432 6239
rect 7380 6196 7432 6205
rect 8852 6196 8904 6248
rect 6920 6128 6972 6180
rect 9404 6196 9456 6248
rect 10048 6196 10100 6248
rect 10324 6196 10376 6248
rect 11888 6196 11940 6248
rect 14004 6239 14056 6248
rect 14004 6205 14013 6239
rect 14013 6205 14047 6239
rect 14047 6205 14056 6239
rect 14004 6196 14056 6205
rect 10968 6128 11020 6180
rect 12348 6171 12400 6180
rect 12348 6137 12357 6171
rect 12357 6137 12391 6171
rect 12391 6137 12400 6171
rect 12348 6128 12400 6137
rect 14188 6128 14240 6180
rect 9956 6060 10008 6112
rect 10048 6103 10100 6112
rect 10048 6069 10057 6103
rect 10057 6069 10091 6103
rect 10091 6069 10100 6103
rect 10048 6060 10100 6069
rect 10416 6103 10468 6112
rect 10416 6069 10425 6103
rect 10425 6069 10459 6103
rect 10459 6069 10468 6103
rect 10416 6060 10468 6069
rect 12808 6103 12860 6112
rect 12808 6069 12817 6103
rect 12817 6069 12851 6103
rect 12851 6069 12860 6103
rect 12808 6060 12860 6069
rect 12992 6060 13044 6112
rect 13820 6060 13872 6112
rect 14096 6103 14148 6112
rect 14096 6069 14105 6103
rect 14105 6069 14139 6103
rect 14139 6069 14148 6103
rect 14096 6060 14148 6069
rect 14832 6060 14884 6112
rect 4100 5958 4152 6010
rect 4164 5958 4216 6010
rect 4228 5958 4280 6010
rect 4292 5958 4344 6010
rect 4356 5958 4408 6010
rect 7802 5958 7854 6010
rect 7866 5958 7918 6010
rect 7930 5958 7982 6010
rect 7994 5958 8046 6010
rect 8058 5958 8110 6010
rect 11504 5958 11556 6010
rect 11568 5958 11620 6010
rect 11632 5958 11684 6010
rect 11696 5958 11748 6010
rect 11760 5958 11812 6010
rect 15206 5958 15258 6010
rect 15270 5958 15322 6010
rect 15334 5958 15386 6010
rect 15398 5958 15450 6010
rect 15462 5958 15514 6010
rect 1124 5899 1176 5908
rect 1124 5865 1133 5899
rect 1133 5865 1167 5899
rect 1167 5865 1176 5899
rect 1124 5856 1176 5865
rect 1860 5856 1912 5908
rect 3700 5856 3752 5908
rect 5632 5899 5684 5908
rect 5632 5865 5641 5899
rect 5641 5865 5675 5899
rect 5675 5865 5684 5899
rect 5632 5856 5684 5865
rect 6828 5856 6880 5908
rect 7104 5899 7156 5908
rect 7104 5865 7113 5899
rect 7113 5865 7147 5899
rect 7147 5865 7156 5899
rect 7104 5856 7156 5865
rect 7196 5856 7248 5908
rect 8944 5856 8996 5908
rect 10048 5856 10100 5908
rect 10692 5856 10744 5908
rect 10968 5899 11020 5908
rect 10968 5865 10977 5899
rect 10977 5865 11011 5899
rect 11011 5865 11020 5899
rect 10968 5856 11020 5865
rect 11888 5856 11940 5908
rect 12256 5856 12308 5908
rect 14832 5856 14884 5908
rect 3240 5831 3292 5840
rect 3240 5797 3249 5831
rect 3249 5797 3283 5831
rect 3283 5797 3292 5831
rect 3240 5788 3292 5797
rect 1308 5763 1360 5772
rect 1308 5729 1317 5763
rect 1317 5729 1351 5763
rect 1351 5729 1360 5763
rect 1308 5720 1360 5729
rect 3516 5763 3568 5772
rect 3516 5729 3525 5763
rect 3525 5729 3559 5763
rect 3559 5729 3568 5763
rect 3516 5720 3568 5729
rect 4620 5720 4672 5772
rect 4896 5652 4948 5704
rect 7656 5720 7708 5772
rect 10324 5788 10376 5840
rect 8576 5720 8628 5772
rect 8852 5720 8904 5772
rect 9312 5720 9364 5772
rect 10876 5788 10928 5840
rect 13820 5788 13872 5840
rect 3056 5584 3108 5636
rect 2964 5516 3016 5568
rect 6736 5652 6788 5704
rect 7472 5652 7524 5704
rect 6736 5516 6788 5568
rect 7564 5559 7616 5568
rect 7564 5525 7573 5559
rect 7573 5525 7607 5559
rect 7607 5525 7616 5559
rect 7564 5516 7616 5525
rect 9404 5652 9456 5704
rect 9496 5652 9548 5704
rect 10232 5695 10284 5704
rect 10232 5661 10241 5695
rect 10241 5661 10275 5695
rect 10275 5661 10284 5695
rect 10232 5652 10284 5661
rect 11336 5763 11388 5772
rect 11336 5729 11345 5763
rect 11345 5729 11379 5763
rect 11379 5729 11388 5763
rect 11336 5720 11388 5729
rect 12716 5720 12768 5772
rect 13544 5720 13596 5772
rect 13912 5763 13964 5772
rect 13912 5729 13921 5763
rect 13921 5729 13955 5763
rect 13955 5729 13964 5763
rect 13912 5720 13964 5729
rect 11152 5652 11204 5704
rect 10140 5584 10192 5636
rect 11980 5652 12032 5704
rect 12532 5652 12584 5704
rect 14004 5695 14056 5704
rect 14004 5661 14013 5695
rect 14013 5661 14047 5695
rect 14047 5661 14056 5695
rect 14004 5652 14056 5661
rect 12624 5584 12676 5636
rect 12900 5584 12952 5636
rect 14556 5695 14608 5704
rect 14556 5661 14565 5695
rect 14565 5661 14599 5695
rect 14599 5661 14608 5695
rect 14556 5652 14608 5661
rect 11244 5516 11296 5568
rect 12256 5516 12308 5568
rect 13728 5516 13780 5568
rect 2249 5414 2301 5466
rect 2313 5414 2365 5466
rect 2377 5414 2429 5466
rect 2441 5414 2493 5466
rect 2505 5414 2557 5466
rect 5951 5414 6003 5466
rect 6015 5414 6067 5466
rect 6079 5414 6131 5466
rect 6143 5414 6195 5466
rect 6207 5414 6259 5466
rect 9653 5414 9705 5466
rect 9717 5414 9769 5466
rect 9781 5414 9833 5466
rect 9845 5414 9897 5466
rect 9909 5414 9961 5466
rect 13355 5414 13407 5466
rect 13419 5414 13471 5466
rect 13483 5414 13535 5466
rect 13547 5414 13599 5466
rect 13611 5414 13663 5466
rect 4712 5312 4764 5364
rect 5172 5312 5224 5364
rect 9312 5312 9364 5364
rect 10600 5312 10652 5364
rect 11152 5312 11204 5364
rect 11520 5312 11572 5364
rect 8852 5244 8904 5296
rect 5448 5219 5500 5228
rect 5448 5185 5457 5219
rect 5457 5185 5491 5219
rect 5491 5185 5500 5219
rect 5448 5176 5500 5185
rect 5632 5176 5684 5228
rect 2136 5015 2188 5024
rect 2136 4981 2145 5015
rect 2145 4981 2179 5015
rect 2179 4981 2188 5015
rect 2136 4972 2188 4981
rect 3056 5151 3108 5160
rect 3056 5117 3065 5151
rect 3065 5117 3099 5151
rect 3099 5117 3108 5151
rect 3056 5108 3108 5117
rect 3700 5108 3752 5160
rect 4712 5108 4764 5160
rect 5172 5151 5224 5160
rect 5172 5117 5181 5151
rect 5181 5117 5215 5151
rect 5215 5117 5224 5151
rect 5172 5108 5224 5117
rect 8944 5176 8996 5228
rect 9496 5176 9548 5228
rect 7564 5108 7616 5160
rect 8576 5108 8628 5160
rect 9128 5108 9180 5160
rect 9404 5108 9456 5160
rect 2688 5040 2740 5092
rect 4252 5040 4304 5092
rect 4436 5040 4488 5092
rect 7288 5040 7340 5092
rect 8208 5040 8260 5092
rect 10140 5040 10192 5092
rect 10232 5083 10284 5092
rect 10232 5049 10241 5083
rect 10241 5049 10275 5083
rect 10275 5049 10284 5083
rect 10232 5040 10284 5049
rect 2964 4972 3016 5024
rect 5264 5015 5316 5024
rect 5264 4981 5273 5015
rect 5273 4981 5307 5015
rect 5307 4981 5316 5015
rect 5264 4972 5316 4981
rect 5540 4972 5592 5024
rect 6184 4972 6236 5024
rect 9496 4972 9548 5024
rect 10324 5015 10376 5024
rect 10324 4981 10333 5015
rect 10333 4981 10367 5015
rect 10367 4981 10376 5015
rect 10324 4972 10376 4981
rect 10508 4972 10560 5024
rect 11060 5176 11112 5228
rect 12348 5312 12400 5364
rect 12532 5312 12584 5364
rect 11428 5108 11480 5160
rect 12624 5176 12676 5228
rect 14096 5176 14148 5228
rect 14924 5176 14976 5228
rect 12164 5108 12216 5160
rect 12256 5108 12308 5160
rect 13728 5108 13780 5160
rect 13912 5108 13964 5160
rect 11060 4972 11112 5024
rect 12256 4972 12308 5024
rect 12348 4972 12400 5024
rect 12716 5015 12768 5024
rect 12716 4981 12725 5015
rect 12725 4981 12759 5015
rect 12759 4981 12768 5015
rect 12716 4972 12768 4981
rect 13084 5015 13136 5024
rect 13084 4981 13093 5015
rect 13093 4981 13127 5015
rect 13127 4981 13136 5015
rect 13084 4972 13136 4981
rect 13912 4972 13964 5024
rect 4100 4870 4152 4922
rect 4164 4870 4216 4922
rect 4228 4870 4280 4922
rect 4292 4870 4344 4922
rect 4356 4870 4408 4922
rect 7802 4870 7854 4922
rect 7866 4870 7918 4922
rect 7930 4870 7982 4922
rect 7994 4870 8046 4922
rect 8058 4870 8110 4922
rect 11504 4870 11556 4922
rect 11568 4870 11620 4922
rect 11632 4870 11684 4922
rect 11696 4870 11748 4922
rect 11760 4870 11812 4922
rect 15206 4870 15258 4922
rect 15270 4870 15322 4922
rect 15334 4870 15386 4922
rect 15398 4870 15450 4922
rect 15462 4870 15514 4922
rect 2136 4768 2188 4820
rect 3884 4811 3936 4820
rect 3884 4777 3893 4811
rect 3893 4777 3927 4811
rect 3927 4777 3936 4811
rect 3884 4768 3936 4777
rect 4620 4768 4672 4820
rect 4896 4811 4948 4820
rect 4896 4777 4905 4811
rect 4905 4777 4939 4811
rect 4939 4777 4948 4811
rect 4896 4768 4948 4777
rect 7380 4811 7432 4820
rect 7380 4777 7389 4811
rect 7389 4777 7423 4811
rect 7423 4777 7432 4811
rect 7380 4768 7432 4777
rect 9036 4768 9088 4820
rect 10048 4768 10100 4820
rect 5264 4700 5316 4752
rect 2504 4607 2556 4616
rect 2504 4573 2513 4607
rect 2513 4573 2547 4607
rect 2547 4573 2556 4607
rect 2504 4564 2556 4573
rect 3700 4564 3752 4616
rect 4344 4607 4396 4616
rect 4344 4573 4353 4607
rect 4353 4573 4387 4607
rect 4387 4573 4396 4607
rect 4344 4564 4396 4573
rect 4436 4607 4488 4616
rect 4436 4573 4445 4607
rect 4445 4573 4479 4607
rect 4479 4573 4488 4607
rect 4436 4564 4488 4573
rect 5448 4564 5500 4616
rect 6184 4675 6236 4684
rect 6184 4641 6193 4675
rect 6193 4641 6227 4675
rect 6227 4641 6236 4675
rect 6184 4632 6236 4641
rect 6828 4632 6880 4684
rect 9036 4675 9088 4684
rect 3516 4496 3568 4548
rect 4252 4496 4304 4548
rect 4528 4496 4580 4548
rect 6184 4496 6236 4548
rect 4896 4428 4948 4480
rect 7012 4428 7064 4480
rect 8208 4564 8260 4616
rect 9036 4641 9054 4675
rect 9054 4641 9088 4675
rect 9036 4632 9088 4641
rect 9128 4675 9180 4684
rect 9128 4641 9137 4675
rect 9137 4641 9171 4675
rect 9171 4641 9180 4675
rect 9128 4632 9180 4641
rect 8668 4564 8720 4616
rect 9956 4564 10008 4616
rect 10600 4700 10652 4752
rect 11244 4768 11296 4820
rect 11520 4768 11572 4820
rect 14188 4768 14240 4820
rect 11428 4700 11480 4752
rect 11244 4632 11296 4684
rect 12072 4700 12124 4752
rect 12624 4632 12676 4684
rect 12900 4632 12952 4684
rect 13176 4675 13228 4684
rect 13176 4641 13185 4675
rect 13185 4641 13219 4675
rect 13219 4641 13228 4675
rect 13176 4632 13228 4641
rect 14372 4632 14424 4684
rect 14648 4632 14700 4684
rect 9496 4496 9548 4548
rect 11520 4564 11572 4616
rect 12164 4564 12216 4616
rect 12256 4564 12308 4616
rect 13084 4564 13136 4616
rect 10784 4496 10836 4548
rect 10048 4428 10100 4480
rect 10876 4428 10928 4480
rect 12072 4428 12124 4480
rect 12808 4471 12860 4480
rect 12808 4437 12817 4471
rect 12817 4437 12851 4471
rect 12851 4437 12860 4471
rect 12808 4428 12860 4437
rect 13084 4428 13136 4480
rect 14464 4607 14516 4616
rect 14464 4573 14473 4607
rect 14473 4573 14507 4607
rect 14507 4573 14516 4607
rect 14464 4564 14516 4573
rect 2249 4326 2301 4378
rect 2313 4326 2365 4378
rect 2377 4326 2429 4378
rect 2441 4326 2493 4378
rect 2505 4326 2557 4378
rect 5951 4326 6003 4378
rect 6015 4326 6067 4378
rect 6079 4326 6131 4378
rect 6143 4326 6195 4378
rect 6207 4326 6259 4378
rect 9653 4326 9705 4378
rect 9717 4326 9769 4378
rect 9781 4326 9833 4378
rect 9845 4326 9897 4378
rect 9909 4326 9961 4378
rect 13355 4326 13407 4378
rect 13419 4326 13471 4378
rect 13483 4326 13535 4378
rect 13547 4326 13599 4378
rect 13611 4326 13663 4378
rect 4344 4224 4396 4276
rect 2688 4088 2740 4140
rect 4252 4131 4304 4140
rect 4252 4097 4261 4131
rect 4261 4097 4295 4131
rect 4295 4097 4304 4131
rect 4252 4088 4304 4097
rect 4436 4088 4488 4140
rect 6736 4156 6788 4208
rect 7012 4156 7064 4208
rect 9404 4224 9456 4276
rect 10140 4224 10192 4276
rect 10876 4224 10928 4276
rect 11520 4224 11572 4276
rect 9128 4199 9180 4208
rect 9128 4165 9137 4199
rect 9137 4165 9171 4199
rect 9171 4165 9180 4199
rect 9128 4156 9180 4165
rect 2596 4020 2648 4072
rect 3240 4020 3292 4072
rect 3976 4020 4028 4072
rect 4068 4063 4120 4072
rect 4068 4029 4077 4063
rect 4077 4029 4111 4063
rect 4111 4029 4120 4063
rect 4068 4020 4120 4029
rect 5724 4020 5776 4072
rect 8760 4088 8812 4140
rect 6184 4020 6236 4072
rect 6644 4020 6696 4072
rect 7196 4063 7248 4072
rect 7196 4029 7205 4063
rect 7205 4029 7239 4063
rect 7239 4029 7248 4063
rect 7196 4020 7248 4029
rect 7472 4063 7524 4072
rect 7472 4029 7481 4063
rect 7481 4029 7515 4063
rect 7515 4029 7524 4063
rect 7472 4020 7524 4029
rect 9128 4020 9180 4072
rect 10048 4131 10100 4140
rect 10048 4097 10057 4131
rect 10057 4097 10091 4131
rect 10091 4097 10100 4131
rect 10048 4088 10100 4097
rect 12164 4088 12216 4140
rect 10232 4063 10284 4072
rect 10232 4029 10241 4063
rect 10241 4029 10275 4063
rect 10275 4029 10284 4063
rect 10232 4020 10284 4029
rect 11060 4020 11112 4072
rect 12532 4088 12584 4140
rect 12716 4088 12768 4140
rect 12808 4088 12860 4140
rect 13084 4131 13136 4140
rect 13084 4097 13093 4131
rect 13093 4097 13127 4131
rect 13127 4097 13136 4131
rect 13084 4088 13136 4097
rect 14096 4131 14148 4140
rect 3424 3884 3476 3936
rect 3884 3927 3936 3936
rect 3884 3893 3893 3927
rect 3893 3893 3927 3927
rect 3927 3893 3936 3927
rect 3884 3884 3936 3893
rect 4896 3927 4948 3936
rect 4896 3893 4905 3927
rect 4905 3893 4939 3927
rect 4939 3893 4948 3927
rect 4896 3884 4948 3893
rect 5356 3927 5408 3936
rect 5356 3893 5365 3927
rect 5365 3893 5399 3927
rect 5399 3893 5408 3927
rect 5356 3884 5408 3893
rect 5448 3927 5500 3936
rect 5448 3893 5457 3927
rect 5457 3893 5491 3927
rect 5491 3893 5500 3927
rect 5448 3884 5500 3893
rect 5816 3927 5868 3936
rect 5816 3893 5825 3927
rect 5825 3893 5859 3927
rect 5859 3893 5868 3927
rect 5816 3884 5868 3893
rect 7196 3884 7248 3936
rect 7472 3884 7524 3936
rect 9220 3927 9272 3936
rect 9220 3893 9229 3927
rect 9229 3893 9263 3927
rect 9263 3893 9272 3927
rect 9220 3884 9272 3893
rect 9404 3884 9456 3936
rect 9772 3884 9824 3936
rect 10968 3927 11020 3936
rect 10968 3893 10977 3927
rect 10977 3893 11011 3927
rect 11011 3893 11020 3927
rect 10968 3884 11020 3893
rect 11060 3927 11112 3936
rect 11060 3893 11069 3927
rect 11069 3893 11103 3927
rect 11103 3893 11112 3927
rect 11060 3884 11112 3893
rect 11888 3952 11940 4004
rect 14096 4097 14105 4131
rect 14105 4097 14139 4131
rect 14139 4097 14148 4131
rect 14096 4088 14148 4097
rect 14648 4088 14700 4140
rect 13912 4063 13964 4072
rect 13912 4029 13921 4063
rect 13921 4029 13955 4063
rect 13955 4029 13964 4063
rect 13912 4020 13964 4029
rect 14004 4020 14056 4072
rect 15108 4020 15160 4072
rect 13360 3952 13412 4004
rect 12164 3927 12216 3936
rect 12164 3893 12173 3927
rect 12173 3893 12207 3927
rect 12207 3893 12216 3927
rect 12164 3884 12216 3893
rect 12256 3884 12308 3936
rect 13176 3884 13228 3936
rect 14556 3884 14608 3936
rect 14832 3884 14884 3936
rect 15108 3884 15160 3936
rect 4100 3782 4152 3834
rect 4164 3782 4216 3834
rect 4228 3782 4280 3834
rect 4292 3782 4344 3834
rect 4356 3782 4408 3834
rect 7802 3782 7854 3834
rect 7866 3782 7918 3834
rect 7930 3782 7982 3834
rect 7994 3782 8046 3834
rect 8058 3782 8110 3834
rect 11504 3782 11556 3834
rect 11568 3782 11620 3834
rect 11632 3782 11684 3834
rect 11696 3782 11748 3834
rect 11760 3782 11812 3834
rect 15206 3782 15258 3834
rect 15270 3782 15322 3834
rect 15334 3782 15386 3834
rect 15398 3782 15450 3834
rect 15462 3782 15514 3834
rect 3608 3680 3660 3732
rect 1124 3544 1176 3596
rect 5816 3680 5868 3732
rect 6644 3680 6696 3732
rect 8852 3723 8904 3732
rect 8852 3689 8861 3723
rect 8861 3689 8895 3723
rect 8895 3689 8904 3723
rect 8852 3680 8904 3689
rect 9864 3680 9916 3732
rect 10048 3680 10100 3732
rect 11152 3680 11204 3732
rect 11796 3680 11848 3732
rect 12992 3680 13044 3732
rect 5080 3612 5132 3664
rect 3976 3544 4028 3596
rect 3056 3476 3108 3528
rect 4344 3476 4396 3528
rect 5356 3544 5408 3596
rect 5448 3544 5500 3596
rect 6184 3612 6236 3664
rect 6736 3612 6788 3664
rect 7380 3612 7432 3664
rect 9680 3612 9732 3664
rect 8760 3587 8812 3596
rect 8760 3553 8769 3587
rect 8769 3553 8803 3587
rect 8803 3553 8812 3587
rect 8760 3544 8812 3553
rect 9588 3587 9640 3596
rect 9588 3553 9597 3587
rect 9597 3553 9631 3587
rect 9631 3553 9640 3587
rect 9588 3544 9640 3553
rect 12532 3655 12584 3664
rect 12532 3621 12541 3655
rect 12541 3621 12575 3655
rect 12575 3621 12584 3655
rect 12532 3612 12584 3621
rect 13084 3612 13136 3664
rect 11888 3544 11940 3596
rect 11980 3587 12032 3596
rect 11980 3553 11989 3587
rect 11989 3553 12023 3587
rect 12023 3553 12032 3587
rect 11980 3544 12032 3553
rect 13176 3587 13228 3596
rect 13176 3553 13185 3587
rect 13185 3553 13219 3587
rect 13219 3553 13228 3587
rect 13176 3544 13228 3553
rect 13912 3680 13964 3732
rect 14096 3587 14148 3596
rect 14096 3553 14105 3587
rect 14105 3553 14139 3587
rect 14139 3553 14148 3587
rect 14096 3544 14148 3553
rect 5540 3476 5592 3528
rect 9772 3408 9824 3460
rect 11244 3476 11296 3528
rect 11152 3408 11204 3460
rect 12164 3408 12216 3460
rect 12256 3408 12308 3460
rect 3148 3340 3200 3392
rect 5816 3340 5868 3392
rect 8392 3383 8444 3392
rect 8392 3349 8401 3383
rect 8401 3349 8435 3383
rect 8435 3349 8444 3383
rect 8392 3340 8444 3349
rect 8484 3340 8536 3392
rect 9680 3340 9732 3392
rect 10968 3340 11020 3392
rect 13176 3340 13228 3392
rect 13360 3340 13412 3392
rect 14188 3340 14240 3392
rect 2249 3238 2301 3290
rect 2313 3238 2365 3290
rect 2377 3238 2429 3290
rect 2441 3238 2493 3290
rect 2505 3238 2557 3290
rect 5951 3238 6003 3290
rect 6015 3238 6067 3290
rect 6079 3238 6131 3290
rect 6143 3238 6195 3290
rect 6207 3238 6259 3290
rect 9653 3238 9705 3290
rect 9717 3238 9769 3290
rect 9781 3238 9833 3290
rect 9845 3238 9897 3290
rect 9909 3238 9961 3290
rect 13355 3238 13407 3290
rect 13419 3238 13471 3290
rect 13483 3238 13535 3290
rect 13547 3238 13599 3290
rect 13611 3238 13663 3290
rect 4988 3179 5040 3188
rect 4988 3145 4997 3179
rect 4997 3145 5031 3179
rect 5031 3145 5040 3179
rect 4988 3136 5040 3145
rect 7380 3136 7432 3188
rect 8852 3136 8904 3188
rect 7012 3068 7064 3120
rect 4344 3043 4396 3052
rect 4344 3009 4353 3043
rect 4353 3009 4387 3043
rect 4387 3009 4396 3043
rect 4344 3000 4396 3009
rect 5724 3000 5776 3052
rect 3240 2932 3292 2984
rect 5816 2975 5868 2984
rect 5816 2941 5825 2975
rect 5825 2941 5859 2975
rect 5859 2941 5868 2975
rect 5816 2932 5868 2941
rect 5908 2975 5960 2984
rect 5908 2941 5917 2975
rect 5917 2941 5951 2975
rect 5951 2941 5960 2975
rect 5908 2932 5960 2941
rect 6736 3000 6788 3052
rect 8484 3000 8536 3052
rect 8944 3000 8996 3052
rect 10232 3136 10284 3188
rect 11980 3136 12032 3188
rect 12900 3136 12952 3188
rect 3792 2796 3844 2848
rect 5080 2864 5132 2916
rect 7564 2864 7616 2916
rect 8484 2864 8536 2916
rect 6552 2839 6604 2848
rect 6552 2805 6561 2839
rect 6561 2805 6595 2839
rect 6595 2805 6604 2839
rect 6552 2796 6604 2805
rect 8760 2975 8812 2984
rect 8760 2941 8769 2975
rect 8769 2941 8803 2975
rect 8803 2941 8812 2975
rect 8760 2932 8812 2941
rect 9588 3043 9640 3052
rect 11060 3068 11112 3120
rect 13176 3068 13228 3120
rect 9588 3009 9622 3043
rect 9622 3009 9640 3043
rect 9588 3000 9640 3009
rect 11336 3000 11388 3052
rect 11796 3000 11848 3052
rect 12256 3000 12308 3052
rect 12440 3043 12492 3052
rect 12440 3009 12449 3043
rect 12449 3009 12483 3043
rect 12483 3009 12492 3043
rect 14648 3111 14700 3120
rect 14648 3077 14657 3111
rect 14657 3077 14691 3111
rect 14691 3077 14700 3111
rect 14648 3068 14700 3077
rect 12440 3000 12492 3009
rect 14096 3043 14148 3052
rect 14096 3009 14105 3043
rect 14105 3009 14139 3043
rect 14139 3009 14148 3043
rect 14096 3000 14148 3009
rect 15568 3000 15620 3052
rect 9772 2975 9824 2984
rect 9772 2941 9781 2975
rect 9781 2941 9815 2975
rect 9815 2941 9824 2975
rect 9772 2932 9824 2941
rect 10876 2975 10928 2984
rect 10876 2941 10885 2975
rect 10885 2941 10919 2975
rect 10919 2941 10928 2975
rect 10876 2932 10928 2941
rect 10968 2932 11020 2984
rect 10232 2796 10284 2848
rect 10784 2796 10836 2848
rect 12532 2975 12584 2984
rect 12532 2941 12566 2975
rect 12566 2941 12584 2975
rect 12532 2932 12584 2941
rect 12716 2975 12768 2984
rect 12716 2941 12725 2975
rect 12725 2941 12759 2975
rect 12759 2941 12768 2975
rect 12716 2932 12768 2941
rect 12256 2796 12308 2848
rect 12716 2796 12768 2848
rect 14648 2864 14700 2916
rect 13820 2796 13872 2848
rect 14188 2796 14240 2848
rect 4100 2694 4152 2746
rect 4164 2694 4216 2746
rect 4228 2694 4280 2746
rect 4292 2694 4344 2746
rect 4356 2694 4408 2746
rect 7802 2694 7854 2746
rect 7866 2694 7918 2746
rect 7930 2694 7982 2746
rect 7994 2694 8046 2746
rect 8058 2694 8110 2746
rect 11504 2694 11556 2746
rect 11568 2694 11620 2746
rect 11632 2694 11684 2746
rect 11696 2694 11748 2746
rect 11760 2694 11812 2746
rect 15206 2694 15258 2746
rect 15270 2694 15322 2746
rect 15334 2694 15386 2746
rect 15398 2694 15450 2746
rect 15462 2694 15514 2746
rect 3056 2592 3108 2644
rect 3148 2592 3200 2644
rect 3148 2499 3200 2508
rect 3148 2465 3166 2499
rect 3166 2465 3200 2499
rect 3148 2456 3200 2465
rect 3240 2499 3292 2508
rect 3240 2465 3249 2499
rect 3249 2465 3283 2499
rect 3283 2465 3292 2499
rect 3240 2456 3292 2465
rect 5908 2592 5960 2644
rect 6552 2567 6604 2576
rect 6552 2533 6561 2567
rect 6561 2533 6595 2567
rect 6595 2533 6604 2567
rect 6552 2524 6604 2533
rect 7748 2524 7800 2576
rect 7288 2456 7340 2508
rect 10876 2592 10928 2644
rect 12716 2592 12768 2644
rect 12992 2592 13044 2644
rect 14096 2592 14148 2644
rect 8300 2567 8352 2576
rect 8300 2533 8309 2567
rect 8309 2533 8343 2567
rect 8343 2533 8352 2567
rect 8300 2524 8352 2533
rect 14556 2567 14608 2576
rect 8484 2456 8536 2508
rect 10600 2456 10652 2508
rect 10692 2499 10744 2508
rect 10692 2465 10701 2499
rect 10701 2465 10735 2499
rect 10735 2465 10744 2499
rect 10692 2456 10744 2465
rect 10968 2456 11020 2508
rect 14556 2533 14565 2567
rect 14565 2533 14599 2567
rect 14599 2533 14608 2567
rect 14556 2524 14608 2533
rect 2964 2431 3016 2440
rect 2964 2397 2973 2431
rect 2973 2397 3007 2431
rect 3007 2397 3016 2431
rect 2964 2388 3016 2397
rect 3884 2388 3936 2440
rect 4160 2431 4212 2440
rect 4160 2397 4169 2431
rect 4169 2397 4203 2431
rect 4203 2397 4212 2431
rect 4160 2388 4212 2397
rect 3700 2320 3752 2372
rect 4160 2252 4212 2304
rect 6736 2252 6788 2304
rect 11428 2456 11480 2508
rect 12532 2456 12584 2508
rect 12992 2456 13044 2508
rect 13084 2388 13136 2440
rect 13268 2456 13320 2508
rect 14372 2456 14424 2508
rect 13820 2431 13872 2440
rect 13820 2397 13829 2431
rect 13829 2397 13863 2431
rect 13863 2397 13872 2431
rect 13820 2388 13872 2397
rect 12900 2320 12952 2372
rect 14464 2320 14516 2372
rect 11520 2252 11572 2304
rect 14188 2295 14240 2304
rect 14188 2261 14197 2295
rect 14197 2261 14231 2295
rect 14231 2261 14240 2295
rect 14188 2252 14240 2261
rect 2249 2150 2301 2202
rect 2313 2150 2365 2202
rect 2377 2150 2429 2202
rect 2441 2150 2493 2202
rect 2505 2150 2557 2202
rect 5951 2150 6003 2202
rect 6015 2150 6067 2202
rect 6079 2150 6131 2202
rect 6143 2150 6195 2202
rect 6207 2150 6259 2202
rect 9653 2150 9705 2202
rect 9717 2150 9769 2202
rect 9781 2150 9833 2202
rect 9845 2150 9897 2202
rect 9909 2150 9961 2202
rect 13355 2150 13407 2202
rect 13419 2150 13471 2202
rect 13483 2150 13535 2202
rect 13547 2150 13599 2202
rect 13611 2150 13663 2202
rect 4896 2048 4948 2100
rect 3240 1912 3292 1964
rect 4160 1844 4212 1896
rect 2964 1776 3016 1828
rect 8668 2048 8720 2100
rect 9496 2048 9548 2100
rect 10692 2048 10744 2100
rect 11520 2048 11572 2100
rect 12808 2091 12860 2100
rect 12808 2057 12817 2091
rect 12817 2057 12851 2091
rect 12851 2057 12860 2091
rect 12808 2048 12860 2057
rect 13176 2048 13228 2100
rect 15568 2048 15620 2100
rect 5632 2023 5684 2032
rect 5632 1989 5641 2023
rect 5641 1989 5675 2023
rect 5675 1989 5684 2023
rect 5632 1980 5684 1989
rect 6368 1980 6420 2032
rect 7196 1980 7248 2032
rect 8760 1980 8812 2032
rect 6092 1955 6144 1964
rect 6092 1921 6101 1955
rect 6101 1921 6135 1955
rect 6135 1921 6144 1955
rect 6092 1912 6144 1921
rect 6828 1912 6880 1964
rect 5264 1887 5316 1896
rect 5264 1853 5282 1887
rect 5282 1853 5316 1887
rect 5264 1844 5316 1853
rect 5356 1887 5408 1896
rect 5356 1853 5365 1887
rect 5365 1853 5399 1887
rect 5399 1853 5408 1887
rect 5356 1844 5408 1853
rect 6184 1844 6236 1896
rect 6736 1844 6788 1896
rect 3240 1751 3292 1760
rect 3240 1717 3249 1751
rect 3249 1717 3283 1751
rect 3283 1717 3292 1751
rect 3240 1708 3292 1717
rect 5264 1708 5316 1760
rect 7748 1708 7800 1760
rect 8484 1887 8536 1896
rect 8484 1853 8493 1887
rect 8493 1853 8527 1887
rect 8527 1853 8536 1887
rect 8484 1844 8536 1853
rect 8668 1844 8720 1896
rect 9220 1844 9272 1896
rect 10140 1912 10192 1964
rect 10232 1912 10284 1964
rect 11152 1912 11204 1964
rect 13084 1980 13136 2032
rect 12440 1912 12492 1964
rect 13360 1980 13412 2032
rect 13636 1980 13688 2032
rect 15016 1980 15068 2032
rect 11244 1844 11296 1896
rect 14188 1844 14240 1896
rect 10048 1776 10100 1828
rect 12440 1776 12492 1828
rect 12716 1819 12768 1828
rect 12716 1785 12725 1819
rect 12725 1785 12759 1819
rect 12759 1785 12768 1819
rect 12716 1776 12768 1785
rect 12992 1776 13044 1828
rect 11428 1708 11480 1760
rect 11888 1708 11940 1760
rect 12072 1708 12124 1760
rect 14004 1708 14056 1760
rect 4100 1606 4152 1658
rect 4164 1606 4216 1658
rect 4228 1606 4280 1658
rect 4292 1606 4344 1658
rect 4356 1606 4408 1658
rect 7802 1606 7854 1658
rect 7866 1606 7918 1658
rect 7930 1606 7982 1658
rect 7994 1606 8046 1658
rect 8058 1606 8110 1658
rect 11504 1606 11556 1658
rect 11568 1606 11620 1658
rect 11632 1606 11684 1658
rect 11696 1606 11748 1658
rect 11760 1606 11812 1658
rect 15206 1606 15258 1658
rect 15270 1606 15322 1658
rect 15334 1606 15386 1658
rect 15398 1606 15450 1658
rect 15462 1606 15514 1658
rect 3148 1504 3200 1556
rect 3792 1547 3844 1556
rect 3792 1513 3801 1547
rect 3801 1513 3835 1547
rect 3835 1513 3844 1547
rect 3792 1504 3844 1513
rect 2780 1411 2832 1420
rect 2780 1377 2789 1411
rect 2789 1377 2823 1411
rect 2823 1377 2832 1411
rect 2780 1368 2832 1377
rect 5264 1504 5316 1556
rect 6276 1504 6328 1556
rect 6920 1504 6972 1556
rect 7472 1504 7524 1556
rect 11888 1504 11940 1556
rect 12716 1504 12768 1556
rect 12808 1504 12860 1556
rect 3240 1300 3292 1352
rect 5356 1436 5408 1488
rect 7564 1436 7616 1488
rect 6092 1368 6144 1420
rect 7196 1368 7248 1420
rect 6184 1300 6236 1352
rect 6644 1343 6696 1352
rect 6644 1309 6653 1343
rect 6653 1309 6687 1343
rect 6687 1309 6696 1343
rect 6644 1300 6696 1309
rect 7012 1300 7064 1352
rect 7472 1343 7524 1352
rect 7472 1309 7481 1343
rect 7481 1309 7515 1343
rect 7515 1309 7524 1343
rect 7472 1300 7524 1309
rect 12256 1436 12308 1488
rect 12992 1479 13044 1488
rect 12992 1445 13001 1479
rect 13001 1445 13035 1479
rect 13035 1445 13044 1479
rect 12992 1436 13044 1445
rect 13268 1504 13320 1556
rect 13728 1504 13780 1556
rect 14372 1547 14424 1556
rect 14372 1513 14381 1547
rect 14381 1513 14415 1547
rect 14415 1513 14424 1547
rect 14372 1504 14424 1513
rect 14648 1547 14700 1556
rect 14648 1513 14657 1547
rect 14657 1513 14691 1547
rect 14691 1513 14700 1547
rect 14648 1504 14700 1513
rect 14740 1504 14792 1556
rect 8668 1368 8720 1420
rect 10508 1411 10560 1420
rect 10508 1377 10517 1411
rect 10517 1377 10551 1411
rect 10551 1377 10560 1411
rect 10508 1368 10560 1377
rect 5724 1232 5776 1284
rect 10600 1343 10652 1352
rect 10600 1309 10609 1343
rect 10609 1309 10643 1343
rect 10643 1309 10652 1343
rect 10600 1300 10652 1309
rect 11428 1300 11480 1352
rect 13084 1343 13136 1352
rect 13084 1309 13093 1343
rect 13093 1309 13127 1343
rect 13127 1309 13136 1343
rect 13084 1300 13136 1309
rect 13176 1300 13228 1352
rect 13912 1275 13964 1284
rect 13912 1241 13921 1275
rect 13921 1241 13955 1275
rect 13955 1241 13964 1275
rect 13912 1232 13964 1241
rect 5632 1207 5684 1216
rect 5632 1173 5641 1207
rect 5641 1173 5675 1207
rect 5675 1173 5684 1207
rect 5632 1164 5684 1173
rect 8392 1164 8444 1216
rect 8484 1207 8536 1216
rect 8484 1173 8493 1207
rect 8493 1173 8527 1207
rect 8527 1173 8536 1207
rect 8484 1164 8536 1173
rect 10140 1207 10192 1216
rect 10140 1173 10149 1207
rect 10149 1173 10183 1207
rect 10183 1173 10192 1207
rect 10140 1164 10192 1173
rect 2249 1062 2301 1114
rect 2313 1062 2365 1114
rect 2377 1062 2429 1114
rect 2441 1062 2493 1114
rect 2505 1062 2557 1114
rect 5951 1062 6003 1114
rect 6015 1062 6067 1114
rect 6079 1062 6131 1114
rect 6143 1062 6195 1114
rect 6207 1062 6259 1114
rect 9653 1062 9705 1114
rect 9717 1062 9769 1114
rect 9781 1062 9833 1114
rect 9845 1062 9897 1114
rect 9909 1062 9961 1114
rect 13355 1062 13407 1114
rect 13419 1062 13471 1114
rect 13483 1062 13535 1114
rect 13547 1062 13599 1114
rect 13611 1062 13663 1114
rect 1124 1003 1176 1012
rect 1124 969 1133 1003
rect 1133 969 1167 1003
rect 1167 969 1176 1003
rect 1124 960 1176 969
rect 3424 1003 3476 1012
rect 3424 969 3433 1003
rect 3433 969 3467 1003
rect 3467 969 3476 1003
rect 3424 960 3476 969
rect 4528 960 4580 1012
rect 5080 960 5132 1012
rect 5632 960 5684 1012
rect 5724 960 5776 1012
rect 6644 960 6696 1012
rect 7196 1003 7248 1012
rect 7196 969 7205 1003
rect 7205 969 7239 1003
rect 7239 969 7248 1003
rect 7196 960 7248 969
rect 7656 960 7708 1012
rect 8484 960 8536 1012
rect 10048 960 10100 1012
rect 10140 960 10192 1012
rect 10324 960 10376 1012
rect 11336 960 11388 1012
rect 12348 960 12400 1012
rect 12440 960 12492 1012
rect 13820 960 13872 1012
rect 14556 960 14608 1012
rect 4712 892 4764 944
rect 2780 824 2832 876
rect 940 799 992 808
rect 940 765 949 799
rect 949 765 983 799
rect 983 765 992 799
rect 940 756 992 765
rect 1952 799 2004 808
rect 1952 765 1961 799
rect 1961 765 1995 799
rect 1995 765 2004 799
rect 1952 756 2004 765
rect 2872 756 2924 808
rect 3976 799 4028 808
rect 3976 765 3985 799
rect 3985 765 4019 799
rect 4019 765 4028 799
rect 3976 756 4028 765
rect 4988 799 5040 808
rect 4988 765 4997 799
rect 4997 765 5031 799
rect 5031 765 5040 799
rect 4988 756 5040 765
rect 6184 756 6236 808
rect 8392 824 8444 876
rect 13912 892 13964 944
rect 7012 799 7064 808
rect 7012 765 7021 799
rect 7021 765 7055 799
rect 7055 765 7064 799
rect 7012 756 7064 765
rect 7380 756 7432 808
rect 7472 756 7524 808
rect 8208 799 8260 808
rect 8208 765 8217 799
rect 8217 765 8251 799
rect 8251 765 8260 799
rect 8208 756 8260 765
rect 8944 688 8996 740
rect 10048 799 10100 808
rect 10048 765 10057 799
rect 10057 765 10091 799
rect 10091 765 10100 799
rect 10048 756 10100 765
rect 10508 756 10560 808
rect 11060 799 11112 808
rect 11060 765 11069 799
rect 11069 765 11103 799
rect 11103 765 11112 799
rect 11060 756 11112 765
rect 12072 799 12124 808
rect 12072 765 12081 799
rect 12081 765 12115 799
rect 12115 765 12124 799
rect 12072 756 12124 765
rect 13084 799 13136 808
rect 13084 765 13093 799
rect 13093 765 13127 799
rect 13127 765 13136 799
rect 13084 756 13136 765
rect 13728 799 13780 808
rect 13728 765 13737 799
rect 13737 765 13771 799
rect 13771 765 13780 799
rect 13728 756 13780 765
rect 14004 756 14056 808
rect 15016 799 15068 808
rect 15016 765 15025 799
rect 15025 765 15059 799
rect 15059 765 15068 799
rect 15016 756 15068 765
rect 14924 688 14976 740
rect 15108 620 15160 672
rect 4100 518 4152 570
rect 4164 518 4216 570
rect 4228 518 4280 570
rect 4292 518 4344 570
rect 4356 518 4408 570
rect 7802 518 7854 570
rect 7866 518 7918 570
rect 7930 518 7982 570
rect 7994 518 8046 570
rect 8058 518 8110 570
rect 11504 518 11556 570
rect 11568 518 11620 570
rect 11632 518 11684 570
rect 11696 518 11748 570
rect 11760 518 11812 570
rect 15206 518 15258 570
rect 15270 518 15322 570
rect 15334 518 15386 570
rect 15398 518 15450 570
rect 15462 518 15514 570
rect 8024 416 8076 468
rect 8208 416 8260 468
<< metal2 >>
rect 754 6800 810 7200
rect 1122 6800 1178 7200
rect 1490 6800 1546 7200
rect 1858 6800 1914 7200
rect 2226 6800 2282 7200
rect 2594 6800 2650 7200
rect 2962 6800 3018 7200
rect 3330 6800 3386 7200
rect 3698 6800 3754 7200
rect 4066 6800 4122 7200
rect 4434 6800 4490 7200
rect 4802 6800 4858 7200
rect 5170 6800 5226 7200
rect 5538 6800 5594 7200
rect 5906 6800 5962 7200
rect 6274 6800 6330 7200
rect 6642 6800 6698 7200
rect 7010 6800 7066 7200
rect 7378 6800 7434 7200
rect 7746 6800 7802 7200
rect 8114 6800 8170 7200
rect 8482 6800 8538 7200
rect 8850 6800 8906 7200
rect 9218 6800 9274 7200
rect 9586 6800 9642 7200
rect 9954 6800 10010 7200
rect 10322 6800 10378 7200
rect 10690 6800 10746 7200
rect 11058 6800 11114 7200
rect 11426 6800 11482 7200
rect 11794 6800 11850 7200
rect 11900 6854 12112 6882
rect 768 6254 796 6800
rect 756 6248 808 6254
rect 756 6190 808 6196
rect 1136 5914 1164 6800
rect 1504 6458 1532 6800
rect 1492 6452 1544 6458
rect 1492 6394 1544 6400
rect 1308 6248 1360 6254
rect 1308 6190 1360 6196
rect 1124 5908 1176 5914
rect 1124 5850 1176 5856
rect 1320 5778 1348 6190
rect 1872 5914 1900 6800
rect 2240 6746 2268 6800
rect 2148 6718 2268 6746
rect 2148 6458 2176 6718
rect 2249 6556 2557 6565
rect 2249 6554 2255 6556
rect 2311 6554 2335 6556
rect 2391 6554 2415 6556
rect 2471 6554 2495 6556
rect 2551 6554 2557 6556
rect 2311 6502 2313 6554
rect 2493 6502 2495 6554
rect 2249 6500 2255 6502
rect 2311 6500 2335 6502
rect 2391 6500 2415 6502
rect 2471 6500 2495 6502
rect 2551 6500 2557 6502
rect 2249 6491 2557 6500
rect 2608 6458 2636 6800
rect 2976 6458 3004 6800
rect 3344 6458 3372 6800
rect 2136 6452 2188 6458
rect 2136 6394 2188 6400
rect 2596 6452 2648 6458
rect 2596 6394 2648 6400
rect 2964 6452 3016 6458
rect 2964 6394 3016 6400
rect 3332 6452 3384 6458
rect 3332 6394 3384 6400
rect 3608 6248 3660 6254
rect 3608 6190 3660 6196
rect 1860 5908 1912 5914
rect 1860 5850 1912 5856
rect 3240 5840 3292 5846
rect 3240 5782 3292 5788
rect 1308 5772 1360 5778
rect 1308 5714 1360 5720
rect 3056 5636 3108 5642
rect 3056 5578 3108 5584
rect 2964 5568 3016 5574
rect 2964 5510 3016 5516
rect 2249 5468 2557 5477
rect 2249 5466 2255 5468
rect 2311 5466 2335 5468
rect 2391 5466 2415 5468
rect 2471 5466 2495 5468
rect 2551 5466 2557 5468
rect 2311 5414 2313 5466
rect 2493 5414 2495 5466
rect 2249 5412 2255 5414
rect 2311 5412 2335 5414
rect 2391 5412 2415 5414
rect 2471 5412 2495 5414
rect 2551 5412 2557 5414
rect 2249 5403 2557 5412
rect 2688 5092 2740 5098
rect 2688 5034 2740 5040
rect 2136 5024 2188 5030
rect 2136 4966 2188 4972
rect 2148 4826 2176 4966
rect 2136 4820 2188 4826
rect 2136 4762 2188 4768
rect 2504 4616 2556 4622
rect 2502 4584 2504 4593
rect 2556 4584 2558 4593
rect 2558 4542 2636 4570
rect 2502 4519 2558 4528
rect 2249 4380 2557 4389
rect 2249 4378 2255 4380
rect 2311 4378 2335 4380
rect 2391 4378 2415 4380
rect 2471 4378 2495 4380
rect 2551 4378 2557 4380
rect 2311 4326 2313 4378
rect 2493 4326 2495 4378
rect 2249 4324 2255 4326
rect 2311 4324 2335 4326
rect 2391 4324 2415 4326
rect 2471 4324 2495 4326
rect 2551 4324 2557 4326
rect 2249 4315 2557 4324
rect 2608 4078 2636 4542
rect 2700 4146 2728 5034
rect 2976 5030 3004 5510
rect 3068 5166 3096 5578
rect 3056 5160 3108 5166
rect 3056 5102 3108 5108
rect 2964 5024 3016 5030
rect 2964 4966 3016 4972
rect 2688 4140 2740 4146
rect 2688 4082 2740 4088
rect 2596 4072 2648 4078
rect 2596 4014 2648 4020
rect 1124 3596 1176 3602
rect 1124 3538 1176 3544
rect 1136 1018 1164 3538
rect 2249 3292 2557 3301
rect 2249 3290 2255 3292
rect 2311 3290 2335 3292
rect 2391 3290 2415 3292
rect 2471 3290 2495 3292
rect 2551 3290 2557 3292
rect 2311 3238 2313 3290
rect 2493 3238 2495 3290
rect 2249 3236 2255 3238
rect 2311 3236 2335 3238
rect 2391 3236 2415 3238
rect 2471 3236 2495 3238
rect 2551 3236 2557 3238
rect 2249 3227 2557 3236
rect 2976 2446 3004 4966
rect 3252 4078 3280 5782
rect 3516 5772 3568 5778
rect 3516 5714 3568 5720
rect 3528 4554 3556 5714
rect 3516 4548 3568 4554
rect 3516 4490 3568 4496
rect 3240 4072 3292 4078
rect 3240 4014 3292 4020
rect 3424 3936 3476 3942
rect 3424 3878 3476 3884
rect 3056 3528 3108 3534
rect 3056 3470 3108 3476
rect 3068 2650 3096 3470
rect 3148 3392 3200 3398
rect 3148 3334 3200 3340
rect 3160 2650 3188 3334
rect 3240 2984 3292 2990
rect 3240 2926 3292 2932
rect 3056 2644 3108 2650
rect 3056 2586 3108 2592
rect 3148 2644 3200 2650
rect 3148 2586 3200 2592
rect 3160 2514 3188 2586
rect 3252 2514 3280 2926
rect 3148 2508 3200 2514
rect 3148 2450 3200 2456
rect 3240 2508 3292 2514
rect 3240 2450 3292 2456
rect 2964 2440 3016 2446
rect 2964 2382 3016 2388
rect 2249 2204 2557 2213
rect 2249 2202 2255 2204
rect 2311 2202 2335 2204
rect 2391 2202 2415 2204
rect 2471 2202 2495 2204
rect 2551 2202 2557 2204
rect 2311 2150 2313 2202
rect 2493 2150 2495 2202
rect 2249 2148 2255 2150
rect 2311 2148 2335 2150
rect 2391 2148 2415 2150
rect 2471 2148 2495 2150
rect 2551 2148 2557 2150
rect 2249 2139 2557 2148
rect 2976 1834 3004 2382
rect 2964 1828 3016 1834
rect 2964 1770 3016 1776
rect 3160 1562 3188 2450
rect 3252 1970 3280 2450
rect 3240 1964 3292 1970
rect 3240 1906 3292 1912
rect 3240 1760 3292 1766
rect 3240 1702 3292 1708
rect 3148 1556 3200 1562
rect 3148 1498 3200 1504
rect 2780 1420 2832 1426
rect 2780 1362 2832 1368
rect 2249 1116 2557 1125
rect 2249 1114 2255 1116
rect 2311 1114 2335 1116
rect 2391 1114 2415 1116
rect 2471 1114 2495 1116
rect 2551 1114 2557 1116
rect 2311 1062 2313 1114
rect 2493 1062 2495 1114
rect 2249 1060 2255 1062
rect 2311 1060 2335 1062
rect 2391 1060 2415 1062
rect 2471 1060 2495 1062
rect 2551 1060 2557 1062
rect 2249 1051 2557 1060
rect 1124 1012 1176 1018
rect 1124 954 1176 960
rect 2792 882 2820 1362
rect 3252 1358 3280 1702
rect 3240 1352 3292 1358
rect 3240 1294 3292 1300
rect 3436 1018 3464 3878
rect 3620 3738 3648 6190
rect 3712 5914 3740 6800
rect 4080 6458 4108 6800
rect 4448 6458 4476 6800
rect 4816 6458 4844 6800
rect 4068 6452 4120 6458
rect 4068 6394 4120 6400
rect 4436 6452 4488 6458
rect 4436 6394 4488 6400
rect 4804 6452 4856 6458
rect 4804 6394 4856 6400
rect 5184 6322 5212 6800
rect 5552 6474 5580 6800
rect 5920 6746 5948 6800
rect 5460 6458 5580 6474
rect 5828 6718 5948 6746
rect 5828 6458 5856 6718
rect 5951 6556 6259 6565
rect 5951 6554 5957 6556
rect 6013 6554 6037 6556
rect 6093 6554 6117 6556
rect 6173 6554 6197 6556
rect 6253 6554 6259 6556
rect 6013 6502 6015 6554
rect 6195 6502 6197 6554
rect 5951 6500 5957 6502
rect 6013 6500 6037 6502
rect 6093 6500 6117 6502
rect 6173 6500 6197 6502
rect 6253 6500 6259 6502
rect 5951 6491 6259 6500
rect 6288 6458 6316 6800
rect 6656 6458 6684 6800
rect 7024 6458 7052 6800
rect 7104 6724 7156 6730
rect 7104 6666 7156 6672
rect 5448 6452 5580 6458
rect 5500 6446 5580 6452
rect 5816 6452 5868 6458
rect 5448 6394 5500 6400
rect 5816 6394 5868 6400
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 6644 6452 6696 6458
rect 6644 6394 6696 6400
rect 7012 6452 7064 6458
rect 7012 6394 7064 6400
rect 5172 6316 5224 6322
rect 5172 6258 5224 6264
rect 3884 6248 3936 6254
rect 3884 6190 3936 6196
rect 4528 6248 4580 6254
rect 4528 6190 4580 6196
rect 4712 6248 4764 6254
rect 4712 6190 4764 6196
rect 5356 6248 5408 6254
rect 5356 6190 5408 6196
rect 6184 6248 6236 6254
rect 6184 6190 6236 6196
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 3700 5908 3752 5914
rect 3700 5850 3752 5856
rect 3700 5160 3752 5166
rect 3700 5102 3752 5108
rect 3712 4622 3740 5102
rect 3896 4826 3924 6190
rect 4100 6012 4408 6021
rect 4100 6010 4106 6012
rect 4162 6010 4186 6012
rect 4242 6010 4266 6012
rect 4322 6010 4346 6012
rect 4402 6010 4408 6012
rect 4162 5958 4164 6010
rect 4344 5958 4346 6010
rect 4100 5956 4106 5958
rect 4162 5956 4186 5958
rect 4242 5956 4266 5958
rect 4322 5956 4346 5958
rect 4402 5956 4408 5958
rect 4100 5947 4408 5956
rect 4252 5092 4304 5098
rect 4436 5092 4488 5098
rect 4304 5052 4436 5080
rect 4252 5034 4304 5040
rect 4436 5034 4488 5040
rect 4100 4924 4408 4933
rect 4100 4922 4106 4924
rect 4162 4922 4186 4924
rect 4242 4922 4266 4924
rect 4322 4922 4346 4924
rect 4402 4922 4408 4924
rect 4162 4870 4164 4922
rect 4344 4870 4346 4922
rect 4100 4868 4106 4870
rect 4162 4868 4186 4870
rect 4242 4868 4266 4870
rect 4322 4868 4346 4870
rect 4402 4868 4408 4870
rect 4100 4859 4408 4868
rect 3884 4820 3936 4826
rect 3884 4762 3936 4768
rect 3700 4616 3752 4622
rect 3700 4558 3752 4564
rect 4344 4616 4396 4622
rect 4344 4558 4396 4564
rect 4436 4616 4488 4622
rect 4436 4558 4488 4564
rect 3608 3732 3660 3738
rect 3608 3674 3660 3680
rect 3712 2378 3740 4558
rect 4252 4548 4304 4554
rect 4252 4490 4304 4496
rect 4264 4146 4292 4490
rect 4356 4282 4384 4558
rect 4344 4276 4396 4282
rect 4344 4218 4396 4224
rect 4448 4146 4476 4558
rect 4540 4554 4568 6190
rect 4620 5772 4672 5778
rect 4620 5714 4672 5720
rect 4632 4826 4660 5714
rect 4724 5370 4752 6190
rect 4988 6180 5040 6186
rect 4988 6122 5040 6128
rect 4896 5704 4948 5710
rect 4896 5646 4948 5652
rect 4712 5364 4764 5370
rect 4712 5306 4764 5312
rect 4712 5160 4764 5166
rect 4712 5102 4764 5108
rect 4620 4820 4672 4826
rect 4620 4762 4672 4768
rect 4528 4548 4580 4554
rect 4528 4490 4580 4496
rect 4632 4434 4660 4762
rect 4540 4406 4660 4434
rect 4252 4140 4304 4146
rect 4252 4082 4304 4088
rect 4436 4140 4488 4146
rect 4436 4082 4488 4088
rect 3976 4072 4028 4078
rect 4068 4072 4120 4078
rect 3976 4014 4028 4020
rect 4066 4040 4068 4049
rect 4120 4040 4122 4049
rect 3884 3936 3936 3942
rect 3884 3878 3936 3884
rect 3792 2848 3844 2854
rect 3792 2790 3844 2796
rect 3700 2372 3752 2378
rect 3700 2314 3752 2320
rect 3712 2281 3740 2314
rect 3698 2272 3754 2281
rect 3698 2207 3754 2216
rect 3804 1562 3832 2790
rect 3896 2446 3924 3878
rect 3988 3602 4016 4014
rect 4066 3975 4122 3984
rect 4100 3836 4408 3845
rect 4100 3834 4106 3836
rect 4162 3834 4186 3836
rect 4242 3834 4266 3836
rect 4322 3834 4346 3836
rect 4402 3834 4408 3836
rect 4162 3782 4164 3834
rect 4344 3782 4346 3834
rect 4100 3780 4106 3782
rect 4162 3780 4186 3782
rect 4242 3780 4266 3782
rect 4322 3780 4346 3782
rect 4402 3780 4408 3782
rect 4100 3771 4408 3780
rect 3976 3596 4028 3602
rect 3976 3538 4028 3544
rect 4344 3528 4396 3534
rect 4448 3516 4476 4082
rect 4396 3488 4476 3516
rect 4344 3470 4396 3476
rect 4356 3058 4384 3470
rect 4344 3052 4396 3058
rect 4344 2994 4396 3000
rect 4100 2748 4408 2757
rect 4100 2746 4106 2748
rect 4162 2746 4186 2748
rect 4242 2746 4266 2748
rect 4322 2746 4346 2748
rect 4402 2746 4408 2748
rect 4162 2694 4164 2746
rect 4344 2694 4346 2746
rect 4100 2692 4106 2694
rect 4162 2692 4186 2694
rect 4242 2692 4266 2694
rect 4322 2692 4346 2694
rect 4402 2692 4408 2694
rect 4100 2683 4408 2692
rect 3884 2440 3936 2446
rect 3884 2382 3936 2388
rect 4160 2440 4212 2446
rect 4160 2382 4212 2388
rect 4172 2310 4200 2382
rect 4160 2304 4212 2310
rect 4160 2246 4212 2252
rect 4172 1902 4200 2246
rect 4160 1896 4212 1902
rect 4160 1838 4212 1844
rect 4100 1660 4408 1669
rect 4100 1658 4106 1660
rect 4162 1658 4186 1660
rect 4242 1658 4266 1660
rect 4322 1658 4346 1660
rect 4402 1658 4408 1660
rect 4162 1606 4164 1658
rect 4344 1606 4346 1658
rect 4100 1604 4106 1606
rect 4162 1604 4186 1606
rect 4242 1604 4266 1606
rect 4322 1604 4346 1606
rect 4402 1604 4408 1606
rect 4100 1595 4408 1604
rect 3792 1556 3844 1562
rect 3792 1498 3844 1504
rect 4540 1018 4568 4406
rect 3424 1012 3476 1018
rect 3424 954 3476 960
rect 4528 1012 4580 1018
rect 4528 954 4580 960
rect 4724 950 4752 5102
rect 4908 4826 4936 5646
rect 4896 4820 4948 4826
rect 4896 4762 4948 4768
rect 4908 4486 4936 4762
rect 4896 4480 4948 4486
rect 4896 4422 4948 4428
rect 4896 3936 4948 3942
rect 4896 3878 4948 3884
rect 4908 2106 4936 3878
rect 5000 3194 5028 6122
rect 5172 5364 5224 5370
rect 5172 5306 5224 5312
rect 5184 5166 5212 5306
rect 5172 5160 5224 5166
rect 5172 5102 5224 5108
rect 5264 5024 5316 5030
rect 5264 4966 5316 4972
rect 5276 4758 5304 4966
rect 5264 4752 5316 4758
rect 5264 4694 5316 4700
rect 5368 3942 5396 6190
rect 5632 5908 5684 5914
rect 5632 5850 5684 5856
rect 5644 5234 5672 5850
rect 6196 5658 6224 6190
rect 6840 5914 6868 6190
rect 6920 6180 6972 6186
rect 6920 6122 6972 6128
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 6736 5704 6788 5710
rect 6196 5630 6316 5658
rect 6736 5646 6788 5652
rect 5951 5468 6259 5477
rect 5951 5466 5957 5468
rect 6013 5466 6037 5468
rect 6093 5466 6117 5468
rect 6173 5466 6197 5468
rect 6253 5466 6259 5468
rect 6013 5414 6015 5466
rect 6195 5414 6197 5466
rect 5951 5412 5957 5414
rect 6013 5412 6037 5414
rect 6093 5412 6117 5414
rect 6173 5412 6197 5414
rect 6253 5412 6259 5414
rect 5951 5403 6259 5412
rect 5448 5228 5500 5234
rect 5448 5170 5500 5176
rect 5632 5228 5684 5234
rect 5632 5170 5684 5176
rect 5460 4622 5488 5170
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 6184 5024 6236 5030
rect 6184 4966 6236 4972
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 5448 3936 5500 3942
rect 5448 3878 5500 3884
rect 5080 3664 5132 3670
rect 5080 3606 5132 3612
rect 4988 3188 5040 3194
rect 4988 3130 5040 3136
rect 5092 2922 5120 3606
rect 5460 3602 5488 3878
rect 5356 3596 5408 3602
rect 5356 3538 5408 3544
rect 5448 3596 5500 3602
rect 5448 3538 5500 3544
rect 5080 2916 5132 2922
rect 5080 2858 5132 2864
rect 4896 2100 4948 2106
rect 4896 2042 4948 2048
rect 5092 1018 5120 2858
rect 5368 2774 5396 3538
rect 5552 3534 5580 4966
rect 6196 4690 6224 4966
rect 6184 4684 6236 4690
rect 6184 4626 6236 4632
rect 6196 4554 6224 4626
rect 6184 4548 6236 4554
rect 6184 4490 6236 4496
rect 5951 4380 6259 4389
rect 5951 4378 5957 4380
rect 6013 4378 6037 4380
rect 6093 4378 6117 4380
rect 6173 4378 6197 4380
rect 6253 4378 6259 4380
rect 6013 4326 6015 4378
rect 6195 4326 6197 4378
rect 5951 4324 5957 4326
rect 6013 4324 6037 4326
rect 6093 4324 6117 4326
rect 6173 4324 6197 4326
rect 6253 4324 6259 4326
rect 5951 4315 6259 4324
rect 5724 4072 5776 4078
rect 5724 4014 5776 4020
rect 6184 4072 6236 4078
rect 6184 4014 6236 4020
rect 5540 3528 5592 3534
rect 5540 3470 5592 3476
rect 5736 3058 5764 4014
rect 5816 3936 5868 3942
rect 5816 3878 5868 3884
rect 5828 3738 5856 3878
rect 5816 3732 5868 3738
rect 5816 3674 5868 3680
rect 6196 3670 6224 4014
rect 6184 3664 6236 3670
rect 6184 3606 6236 3612
rect 5816 3392 5868 3398
rect 5816 3334 5868 3340
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 5828 2990 5856 3334
rect 5951 3292 6259 3301
rect 5951 3290 5957 3292
rect 6013 3290 6037 3292
rect 6093 3290 6117 3292
rect 6173 3290 6197 3292
rect 6253 3290 6259 3292
rect 6013 3238 6015 3290
rect 6195 3238 6197 3290
rect 5951 3236 5957 3238
rect 6013 3236 6037 3238
rect 6093 3236 6117 3238
rect 6173 3236 6197 3238
rect 6253 3236 6259 3238
rect 5951 3227 6259 3236
rect 5816 2984 5868 2990
rect 5816 2926 5868 2932
rect 5908 2984 5960 2990
rect 5908 2926 5960 2932
rect 5920 2774 5948 2926
rect 5368 2746 5948 2774
rect 5368 1902 5396 2746
rect 5920 2650 5948 2746
rect 5908 2644 5960 2650
rect 5908 2586 5960 2592
rect 5630 2272 5686 2281
rect 5630 2207 5686 2216
rect 5644 2038 5672 2207
rect 5951 2204 6259 2213
rect 5951 2202 5957 2204
rect 6013 2202 6037 2204
rect 6093 2202 6117 2204
rect 6173 2202 6197 2204
rect 6253 2202 6259 2204
rect 6013 2150 6015 2202
rect 6195 2150 6197 2202
rect 5951 2148 5957 2150
rect 6013 2148 6037 2150
rect 6093 2148 6117 2150
rect 6173 2148 6197 2150
rect 6253 2148 6259 2150
rect 5951 2139 6259 2148
rect 5632 2032 5684 2038
rect 5632 1974 5684 1980
rect 6092 1964 6144 1970
rect 6092 1906 6144 1912
rect 5264 1896 5316 1902
rect 5264 1838 5316 1844
rect 5356 1896 5408 1902
rect 5356 1838 5408 1844
rect 5276 1766 5304 1838
rect 5264 1760 5316 1766
rect 5264 1702 5316 1708
rect 5276 1562 5304 1702
rect 5264 1556 5316 1562
rect 5264 1498 5316 1504
rect 5368 1494 5396 1838
rect 5356 1488 5408 1494
rect 5356 1430 5408 1436
rect 6104 1426 6132 1906
rect 6184 1896 6236 1902
rect 6184 1838 6236 1844
rect 6092 1420 6144 1426
rect 6092 1362 6144 1368
rect 6196 1358 6224 1838
rect 6288 1562 6316 5630
rect 6748 5574 6776 5646
rect 6736 5568 6788 5574
rect 6736 5510 6788 5516
rect 6366 4720 6422 4729
rect 6366 4655 6422 4664
rect 6380 2038 6408 4655
rect 6748 4214 6776 5510
rect 6828 4684 6880 4690
rect 6828 4626 6880 4632
rect 6736 4208 6788 4214
rect 6736 4150 6788 4156
rect 6644 4072 6696 4078
rect 6644 4014 6696 4020
rect 6656 3738 6684 4014
rect 6644 3732 6696 3738
rect 6644 3674 6696 3680
rect 6736 3664 6788 3670
rect 6840 3641 6868 4626
rect 6736 3606 6788 3612
rect 6826 3632 6882 3641
rect 6748 3058 6776 3606
rect 6826 3567 6882 3576
rect 6736 3052 6788 3058
rect 6736 2994 6788 3000
rect 6552 2848 6604 2854
rect 6552 2790 6604 2796
rect 6564 2582 6592 2790
rect 6552 2576 6604 2582
rect 6552 2518 6604 2524
rect 6736 2304 6788 2310
rect 6736 2246 6788 2252
rect 6368 2032 6420 2038
rect 6368 1974 6420 1980
rect 6748 1902 6776 2246
rect 6826 2000 6882 2009
rect 6826 1935 6828 1944
rect 6880 1935 6882 1944
rect 6828 1906 6880 1912
rect 6736 1896 6788 1902
rect 6736 1838 6788 1844
rect 6932 1562 6960 6122
rect 7116 5914 7144 6666
rect 7392 6458 7420 6800
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 7380 6452 7432 6458
rect 7380 6394 7432 6400
rect 7380 6248 7432 6254
rect 7380 6190 7432 6196
rect 7104 5908 7156 5914
rect 7104 5850 7156 5856
rect 7196 5908 7248 5914
rect 7196 5850 7248 5856
rect 7208 4978 7236 5850
rect 7288 5092 7340 5098
rect 7288 5034 7340 5040
rect 7116 4950 7236 4978
rect 7116 4604 7144 4950
rect 7116 4576 7236 4604
rect 7012 4480 7064 4486
rect 7064 4440 7144 4468
rect 7012 4422 7064 4428
rect 7012 4208 7064 4214
rect 7012 4150 7064 4156
rect 7024 3126 7052 4150
rect 7012 3120 7064 3126
rect 7012 3062 7064 3068
rect 7116 2774 7144 4440
rect 7208 4078 7236 4576
rect 7196 4072 7248 4078
rect 7196 4014 7248 4020
rect 7208 3942 7236 4014
rect 7196 3936 7248 3942
rect 7196 3878 7248 3884
rect 7024 2746 7144 2774
rect 6276 1556 6328 1562
rect 6276 1498 6328 1504
rect 6920 1556 6972 1562
rect 6920 1498 6972 1504
rect 7024 1358 7052 2746
rect 7300 2514 7328 5034
rect 7392 4826 7420 6190
rect 7484 5710 7512 6734
rect 7760 6458 7788 6800
rect 8128 6662 8156 6800
rect 8116 6656 8168 6662
rect 8116 6598 8168 6604
rect 7748 6452 7800 6458
rect 7748 6394 7800 6400
rect 8496 6322 8524 6800
rect 8864 6390 8892 6800
rect 8852 6384 8904 6390
rect 8852 6326 8904 6332
rect 8944 6384 8996 6390
rect 8944 6326 8996 6332
rect 8484 6316 8536 6322
rect 8484 6258 8536 6264
rect 8852 6248 8904 6254
rect 8852 6190 8904 6196
rect 7802 6012 8110 6021
rect 7802 6010 7808 6012
rect 7864 6010 7888 6012
rect 7944 6010 7968 6012
rect 8024 6010 8048 6012
rect 8104 6010 8110 6012
rect 7864 5958 7866 6010
rect 8046 5958 8048 6010
rect 7802 5956 7808 5958
rect 7864 5956 7888 5958
rect 7944 5956 7968 5958
rect 8024 5956 8048 5958
rect 8104 5956 8110 5958
rect 7802 5947 8110 5956
rect 8864 5778 8892 6190
rect 8956 5914 8984 6326
rect 8944 5908 8996 5914
rect 8944 5850 8996 5856
rect 7656 5772 7708 5778
rect 7656 5714 7708 5720
rect 8576 5772 8628 5778
rect 8576 5714 8628 5720
rect 8852 5772 8904 5778
rect 8852 5714 8904 5720
rect 7472 5704 7524 5710
rect 7472 5646 7524 5652
rect 7564 5568 7616 5574
rect 7564 5510 7616 5516
rect 7576 5166 7604 5510
rect 7564 5160 7616 5166
rect 7564 5102 7616 5108
rect 7380 4820 7432 4826
rect 7380 4762 7432 4768
rect 7472 4072 7524 4078
rect 7392 4032 7472 4060
rect 7392 3670 7420 4032
rect 7472 4014 7524 4020
rect 7472 3936 7524 3942
rect 7472 3878 7524 3884
rect 7380 3664 7432 3670
rect 7380 3606 7432 3612
rect 7392 3194 7420 3606
rect 7380 3188 7432 3194
rect 7380 3130 7432 3136
rect 7288 2508 7340 2514
rect 7288 2450 7340 2456
rect 7196 2032 7248 2038
rect 7196 1974 7248 1980
rect 7208 1426 7236 1974
rect 7484 1562 7512 3878
rect 7564 2916 7616 2922
rect 7564 2858 7616 2864
rect 7472 1556 7524 1562
rect 7392 1516 7472 1544
rect 7196 1420 7248 1426
rect 7196 1362 7248 1368
rect 6184 1352 6236 1358
rect 6184 1294 6236 1300
rect 6644 1352 6696 1358
rect 6644 1294 6696 1300
rect 7012 1352 7064 1358
rect 7012 1294 7064 1300
rect 5724 1284 5776 1290
rect 5724 1226 5776 1232
rect 5632 1216 5684 1222
rect 5632 1158 5684 1164
rect 5644 1018 5672 1158
rect 5736 1018 5764 1226
rect 5951 1116 6259 1125
rect 5951 1114 5957 1116
rect 6013 1114 6037 1116
rect 6093 1114 6117 1116
rect 6173 1114 6197 1116
rect 6253 1114 6259 1116
rect 6013 1062 6015 1114
rect 6195 1062 6197 1114
rect 5951 1060 5957 1062
rect 6013 1060 6037 1062
rect 6093 1060 6117 1062
rect 6173 1060 6197 1062
rect 6253 1060 6259 1062
rect 5951 1051 6259 1060
rect 6656 1018 6684 1294
rect 7208 1018 7236 1362
rect 5080 1012 5132 1018
rect 5080 954 5132 960
rect 5632 1012 5684 1018
rect 5632 954 5684 960
rect 5724 1012 5776 1018
rect 5724 954 5776 960
rect 6644 1012 6696 1018
rect 6644 954 6696 960
rect 7196 1012 7248 1018
rect 7196 954 7248 960
rect 4712 944 4764 950
rect 4712 886 4764 892
rect 2780 876 2832 882
rect 2780 818 2832 824
rect 7392 814 7420 1516
rect 7472 1498 7524 1504
rect 7576 1494 7604 2858
rect 7564 1488 7616 1494
rect 7564 1430 7616 1436
rect 7472 1352 7524 1358
rect 7472 1294 7524 1300
rect 7484 814 7512 1294
rect 7668 1018 7696 5714
rect 8588 5166 8616 5714
rect 8852 5296 8904 5302
rect 8852 5238 8904 5244
rect 8576 5160 8628 5166
rect 8576 5102 8628 5108
rect 8208 5092 8260 5098
rect 8208 5034 8260 5040
rect 7802 4924 8110 4933
rect 7802 4922 7808 4924
rect 7864 4922 7888 4924
rect 7944 4922 7968 4924
rect 8024 4922 8048 4924
rect 8104 4922 8110 4924
rect 7864 4870 7866 4922
rect 8046 4870 8048 4922
rect 7802 4868 7808 4870
rect 7864 4868 7888 4870
rect 7944 4868 7968 4870
rect 8024 4868 8048 4870
rect 8104 4868 8110 4870
rect 7802 4859 8110 4868
rect 8220 4622 8248 5034
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 7802 3836 8110 3845
rect 7802 3834 7808 3836
rect 7864 3834 7888 3836
rect 7944 3834 7968 3836
rect 8024 3834 8048 3836
rect 8104 3834 8110 3836
rect 7864 3782 7866 3834
rect 8046 3782 8048 3834
rect 7802 3780 7808 3782
rect 7864 3780 7888 3782
rect 7944 3780 7968 3782
rect 8024 3780 8048 3782
rect 8104 3780 8110 3782
rect 7802 3771 8110 3780
rect 8392 3392 8444 3398
rect 8392 3334 8444 3340
rect 8484 3392 8536 3398
rect 8484 3334 8536 3340
rect 8404 2774 8432 3334
rect 8496 3058 8524 3334
rect 8484 3052 8536 3058
rect 8484 2994 8536 3000
rect 8484 2916 8536 2922
rect 8588 2904 8616 5102
rect 8668 4616 8720 4622
rect 8668 4558 8720 4564
rect 8536 2876 8616 2904
rect 8484 2858 8536 2864
rect 7802 2748 8110 2757
rect 7802 2746 7808 2748
rect 7864 2746 7888 2748
rect 7944 2746 7968 2748
rect 8024 2746 8048 2748
rect 8104 2746 8110 2748
rect 7864 2694 7866 2746
rect 8046 2694 8048 2746
rect 7802 2692 7808 2694
rect 7864 2692 7888 2694
rect 7944 2692 7968 2694
rect 8024 2692 8048 2694
rect 8104 2692 8110 2694
rect 7802 2683 8110 2692
rect 8312 2746 8432 2774
rect 8312 2582 8340 2746
rect 7748 2576 7800 2582
rect 7748 2518 7800 2524
rect 8300 2576 8352 2582
rect 8300 2518 8352 2524
rect 7760 1766 7788 2518
rect 8484 2508 8536 2514
rect 8484 2450 8536 2456
rect 8496 1902 8524 2450
rect 8680 2417 8708 4558
rect 8758 4176 8814 4185
rect 8758 4111 8760 4120
rect 8812 4111 8814 4120
rect 8760 4082 8812 4088
rect 8864 3738 8892 5238
rect 8944 5228 8996 5234
rect 8944 5170 8996 5176
rect 8852 3732 8904 3738
rect 8852 3674 8904 3680
rect 8760 3596 8812 3602
rect 8760 3538 8812 3544
rect 8772 3097 8800 3538
rect 8864 3194 8892 3674
rect 8852 3188 8904 3194
rect 8852 3130 8904 3136
rect 8758 3088 8814 3097
rect 8956 3058 8984 5170
rect 9128 5160 9180 5166
rect 9128 5102 9180 5108
rect 9036 4820 9088 4826
rect 9036 4762 9088 4768
rect 9048 4690 9076 4762
rect 9140 4690 9168 5102
rect 9036 4684 9088 4690
rect 9036 4626 9088 4632
rect 9128 4684 9180 4690
rect 9128 4626 9180 4632
rect 9048 3924 9076 4626
rect 9128 4208 9180 4214
rect 9128 4150 9180 4156
rect 9140 4078 9168 4150
rect 9128 4072 9180 4078
rect 9232 4049 9260 6800
rect 9600 6610 9628 6800
rect 9968 6746 9996 6800
rect 9968 6718 10088 6746
rect 9416 6582 9628 6610
rect 9416 6254 9444 6582
rect 9653 6556 9961 6565
rect 9653 6554 9659 6556
rect 9715 6554 9739 6556
rect 9795 6554 9819 6556
rect 9875 6554 9899 6556
rect 9955 6554 9961 6556
rect 9715 6502 9717 6554
rect 9897 6502 9899 6554
rect 9653 6500 9659 6502
rect 9715 6500 9739 6502
rect 9795 6500 9819 6502
rect 9875 6500 9899 6502
rect 9955 6500 9961 6502
rect 9653 6491 9961 6500
rect 10060 6254 10088 6718
rect 10336 6254 10364 6800
rect 9404 6248 9456 6254
rect 9404 6190 9456 6196
rect 10048 6248 10100 6254
rect 10048 6190 10100 6196
rect 10324 6248 10376 6254
rect 10324 6190 10376 6196
rect 9956 6112 10008 6118
rect 9956 6054 10008 6060
rect 10048 6112 10100 6118
rect 10048 6054 10100 6060
rect 10416 6112 10468 6118
rect 10416 6054 10468 6060
rect 9312 5772 9364 5778
rect 9312 5714 9364 5720
rect 9324 5370 9352 5714
rect 9404 5704 9456 5710
rect 9404 5646 9456 5652
rect 9496 5704 9548 5710
rect 9496 5646 9548 5652
rect 9968 5658 9996 6054
rect 10060 5914 10088 6054
rect 10048 5908 10100 5914
rect 10048 5850 10100 5856
rect 10324 5840 10376 5846
rect 10324 5782 10376 5788
rect 10232 5704 10284 5710
rect 9312 5364 9364 5370
rect 9312 5306 9364 5312
rect 9416 5166 9444 5646
rect 9508 5234 9536 5646
rect 9968 5630 10088 5658
rect 10232 5646 10284 5652
rect 9653 5468 9961 5477
rect 9653 5466 9659 5468
rect 9715 5466 9739 5468
rect 9795 5466 9819 5468
rect 9875 5466 9899 5468
rect 9955 5466 9961 5468
rect 9715 5414 9717 5466
rect 9897 5414 9899 5466
rect 9653 5412 9659 5414
rect 9715 5412 9739 5414
rect 9795 5412 9819 5414
rect 9875 5412 9899 5414
rect 9955 5412 9961 5414
rect 9653 5403 9961 5412
rect 9496 5228 9548 5234
rect 9496 5170 9548 5176
rect 9404 5160 9456 5166
rect 9404 5102 9456 5108
rect 9416 4282 9444 5102
rect 9496 5024 9548 5030
rect 9496 4966 9548 4972
rect 9508 4554 9536 4966
rect 10060 4826 10088 5630
rect 10140 5636 10192 5642
rect 10140 5578 10192 5584
rect 10152 5098 10180 5578
rect 10244 5098 10272 5646
rect 10140 5092 10192 5098
rect 10140 5034 10192 5040
rect 10232 5092 10284 5098
rect 10232 5034 10284 5040
rect 10336 5030 10364 5782
rect 10324 5024 10376 5030
rect 10324 4966 10376 4972
rect 10048 4820 10100 4826
rect 10048 4762 10100 4768
rect 10046 4720 10102 4729
rect 9968 4678 10046 4706
rect 9968 4622 9996 4678
rect 10046 4655 10102 4664
rect 9956 4616 10008 4622
rect 9956 4558 10008 4564
rect 9496 4548 9548 4554
rect 9496 4490 9548 4496
rect 10048 4480 10100 4486
rect 10048 4422 10100 4428
rect 9653 4380 9961 4389
rect 9653 4378 9659 4380
rect 9715 4378 9739 4380
rect 9795 4378 9819 4380
rect 9875 4378 9899 4380
rect 9955 4378 9961 4380
rect 9715 4326 9717 4378
rect 9897 4326 9899 4378
rect 9653 4324 9659 4326
rect 9715 4324 9739 4326
rect 9795 4324 9819 4326
rect 9875 4324 9899 4326
rect 9955 4324 9961 4326
rect 9653 4315 9961 4324
rect 9404 4276 9456 4282
rect 10060 4264 10088 4422
rect 9404 4218 9456 4224
rect 9968 4236 10088 4264
rect 10140 4276 10192 4282
rect 9402 4176 9458 4185
rect 9402 4111 9458 4120
rect 9128 4014 9180 4020
rect 9218 4040 9274 4049
rect 9218 3975 9274 3984
rect 9416 3942 9444 4111
rect 9220 3936 9272 3942
rect 9048 3896 9220 3924
rect 9220 3878 9272 3884
rect 9404 3936 9456 3942
rect 9772 3936 9824 3942
rect 9404 3878 9456 3884
rect 9692 3896 9772 3924
rect 8758 3023 8814 3032
rect 8944 3052 8996 3058
rect 8944 2994 8996 3000
rect 8760 2984 8812 2990
rect 8760 2926 8812 2932
rect 8666 2408 8722 2417
rect 8666 2343 8722 2352
rect 8680 2106 8708 2343
rect 8668 2100 8720 2106
rect 8668 2042 8720 2048
rect 8772 2038 8800 2926
rect 8760 2032 8812 2038
rect 8760 1974 8812 1980
rect 9232 1902 9260 3878
rect 9692 3670 9720 3896
rect 9772 3878 9824 3884
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 9680 3664 9732 3670
rect 9680 3606 9732 3612
rect 9588 3596 9640 3602
rect 9588 3538 9640 3544
rect 9600 3346 9628 3538
rect 9678 3496 9734 3505
rect 9876 3482 9904 3674
rect 9784 3466 9904 3482
rect 9678 3431 9734 3440
rect 9772 3460 9904 3466
rect 9692 3398 9720 3431
rect 9824 3454 9904 3460
rect 9968 3482 9996 4236
rect 10140 4218 10192 4224
rect 10048 4140 10100 4146
rect 10048 4082 10100 4088
rect 10060 3738 10088 4082
rect 10048 3732 10100 3738
rect 10048 3674 10100 3680
rect 9968 3454 10088 3482
rect 9772 3402 9824 3408
rect 9508 3318 9628 3346
rect 9680 3392 9732 3398
rect 9680 3334 9732 3340
rect 9508 2938 9536 3318
rect 9653 3292 9961 3301
rect 9653 3290 9659 3292
rect 9715 3290 9739 3292
rect 9795 3290 9819 3292
rect 9875 3290 9899 3292
rect 9955 3290 9961 3292
rect 9715 3238 9717 3290
rect 9897 3238 9899 3290
rect 9653 3236 9659 3238
rect 9715 3236 9739 3238
rect 9795 3236 9819 3238
rect 9875 3236 9899 3238
rect 9955 3236 9961 3238
rect 9653 3227 9961 3236
rect 9586 3088 9642 3097
rect 9586 3023 9588 3032
rect 9640 3023 9642 3032
rect 9588 2994 9640 3000
rect 9772 2984 9824 2990
rect 9508 2932 9772 2938
rect 9508 2926 9824 2932
rect 9508 2910 9812 2926
rect 9508 2106 9536 2910
rect 9653 2204 9961 2213
rect 9653 2202 9659 2204
rect 9715 2202 9739 2204
rect 9795 2202 9819 2204
rect 9875 2202 9899 2204
rect 9955 2202 9961 2204
rect 9715 2150 9717 2202
rect 9897 2150 9899 2202
rect 9653 2148 9659 2150
rect 9715 2148 9739 2150
rect 9795 2148 9819 2150
rect 9875 2148 9899 2150
rect 9955 2148 9961 2150
rect 9653 2139 9961 2148
rect 9496 2100 9548 2106
rect 9496 2042 9548 2048
rect 8484 1896 8536 1902
rect 8484 1838 8536 1844
rect 8668 1896 8720 1902
rect 8668 1838 8720 1844
rect 9220 1896 9272 1902
rect 9220 1838 9272 1844
rect 7748 1760 7800 1766
rect 7748 1702 7800 1708
rect 7802 1660 8110 1669
rect 7802 1658 7808 1660
rect 7864 1658 7888 1660
rect 7944 1658 7968 1660
rect 8024 1658 8048 1660
rect 8104 1658 8110 1660
rect 7864 1606 7866 1658
rect 8046 1606 8048 1658
rect 7802 1604 7808 1606
rect 7864 1604 7888 1606
rect 7944 1604 7968 1606
rect 8024 1604 8048 1606
rect 8104 1604 8110 1606
rect 7802 1595 8110 1604
rect 8680 1426 8708 1838
rect 10060 1834 10088 3454
rect 10152 1970 10180 4218
rect 10232 4072 10284 4078
rect 10232 4014 10284 4020
rect 10244 3194 10272 4014
rect 10232 3188 10284 3194
rect 10232 3130 10284 3136
rect 10232 2848 10284 2854
rect 10232 2790 10284 2796
rect 10244 1970 10272 2790
rect 10140 1964 10192 1970
rect 10140 1906 10192 1912
rect 10232 1964 10284 1970
rect 10232 1906 10284 1912
rect 10048 1828 10100 1834
rect 10048 1770 10100 1776
rect 8668 1420 8720 1426
rect 8668 1362 8720 1368
rect 8392 1216 8444 1222
rect 8392 1158 8444 1164
rect 8484 1216 8536 1222
rect 8484 1158 8536 1164
rect 7656 1012 7708 1018
rect 7656 954 7708 960
rect 8404 882 8432 1158
rect 8496 1018 8524 1158
rect 9653 1116 9961 1125
rect 9653 1114 9659 1116
rect 9715 1114 9739 1116
rect 9795 1114 9819 1116
rect 9875 1114 9899 1116
rect 9955 1114 9961 1116
rect 9715 1062 9717 1114
rect 9897 1062 9899 1114
rect 9653 1060 9659 1062
rect 9715 1060 9739 1062
rect 9795 1060 9819 1062
rect 9875 1060 9899 1062
rect 9955 1060 9961 1062
rect 9653 1051 9961 1060
rect 10060 1018 10088 1770
rect 10140 1216 10192 1222
rect 10140 1158 10192 1164
rect 10152 1018 10180 1158
rect 10336 1018 10364 4966
rect 10428 3505 10456 6054
rect 10704 5914 10732 6800
rect 10876 6792 10928 6798
rect 10876 6734 10928 6740
rect 10692 5908 10744 5914
rect 10692 5850 10744 5856
rect 10888 5846 10916 6734
rect 10968 6180 11020 6186
rect 10968 6122 11020 6128
rect 10980 5914 11008 6122
rect 10968 5908 11020 5914
rect 10968 5850 11020 5856
rect 10876 5840 10928 5846
rect 10876 5782 10928 5788
rect 10600 5364 10652 5370
rect 10600 5306 10652 5312
rect 10508 5024 10560 5030
rect 10508 4966 10560 4972
rect 10414 3496 10470 3505
rect 10414 3431 10470 3440
rect 10520 3097 10548 4966
rect 10612 4758 10640 5306
rect 11072 5234 11100 6800
rect 11440 5794 11468 6800
rect 11808 6746 11836 6800
rect 11900 6746 11928 6854
rect 11808 6718 11928 6746
rect 11980 6656 12032 6662
rect 11980 6598 12032 6604
rect 11992 6458 12020 6598
rect 11980 6452 12032 6458
rect 11980 6394 12032 6400
rect 11888 6248 11940 6254
rect 11888 6190 11940 6196
rect 11504 6012 11812 6021
rect 11504 6010 11510 6012
rect 11566 6010 11590 6012
rect 11646 6010 11670 6012
rect 11726 6010 11750 6012
rect 11806 6010 11812 6012
rect 11566 5958 11568 6010
rect 11748 5958 11750 6010
rect 11504 5956 11510 5958
rect 11566 5956 11590 5958
rect 11646 5956 11670 5958
rect 11726 5956 11750 5958
rect 11806 5956 11812 5958
rect 11504 5947 11812 5956
rect 11900 5914 11928 6190
rect 11888 5908 11940 5914
rect 11888 5850 11940 5856
rect 11336 5772 11388 5778
rect 11440 5766 11560 5794
rect 11336 5714 11388 5720
rect 11152 5704 11204 5710
rect 11152 5646 11204 5652
rect 11164 5370 11192 5646
rect 11244 5568 11296 5574
rect 11244 5510 11296 5516
rect 11152 5364 11204 5370
rect 11152 5306 11204 5312
rect 11060 5228 11112 5234
rect 11060 5170 11112 5176
rect 11060 5024 11112 5030
rect 11060 4966 11112 4972
rect 10600 4752 10652 4758
rect 10600 4694 10652 4700
rect 10506 3088 10562 3097
rect 10506 3023 10562 3032
rect 10612 2514 10640 4694
rect 10784 4548 10836 4554
rect 10784 4490 10836 4496
rect 10796 2854 10824 4490
rect 10876 4480 10928 4486
rect 10876 4422 10928 4428
rect 10888 4282 10916 4422
rect 10876 4276 10928 4282
rect 10876 4218 10928 4224
rect 11072 4078 11100 4966
rect 11060 4072 11112 4078
rect 11060 4014 11112 4020
rect 10968 3936 11020 3942
rect 10968 3878 11020 3884
rect 11060 3936 11112 3942
rect 11060 3878 11112 3884
rect 10980 3398 11008 3878
rect 10968 3392 11020 3398
rect 10968 3334 11020 3340
rect 11072 3126 11100 3878
rect 11164 3738 11192 5306
rect 11256 4826 11284 5510
rect 11244 4820 11296 4826
rect 11244 4762 11296 4768
rect 11244 4684 11296 4690
rect 11244 4626 11296 4632
rect 11256 3913 11284 4626
rect 11242 3904 11298 3913
rect 11242 3839 11298 3848
rect 11152 3732 11204 3738
rect 11152 3674 11204 3680
rect 11256 3534 11284 3839
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 11152 3460 11204 3466
rect 11152 3402 11204 3408
rect 11060 3120 11112 3126
rect 11060 3062 11112 3068
rect 10876 2984 10928 2990
rect 10876 2926 10928 2932
rect 10968 2984 11020 2990
rect 10968 2926 11020 2932
rect 10784 2848 10836 2854
rect 10784 2790 10836 2796
rect 10888 2650 10916 2926
rect 10876 2644 10928 2650
rect 10876 2586 10928 2592
rect 10980 2514 11008 2926
rect 10600 2508 10652 2514
rect 10600 2450 10652 2456
rect 10692 2508 10744 2514
rect 10692 2450 10744 2456
rect 10968 2508 11020 2514
rect 10968 2450 11020 2456
rect 10508 1420 10560 1426
rect 10508 1362 10560 1368
rect 8484 1012 8536 1018
rect 8484 954 8536 960
rect 10048 1012 10100 1018
rect 10048 954 10100 960
rect 10140 1012 10192 1018
rect 10140 954 10192 960
rect 10324 1012 10376 1018
rect 10324 954 10376 960
rect 8392 876 8444 882
rect 8392 818 8444 824
rect 10520 814 10548 1362
rect 10612 1358 10640 2450
rect 10704 2106 10732 2450
rect 10692 2100 10744 2106
rect 10692 2042 10744 2048
rect 11164 1970 11192 3402
rect 11152 1964 11204 1970
rect 11152 1906 11204 1912
rect 11256 1902 11284 3470
rect 11348 3058 11376 5714
rect 11532 5370 11560 5766
rect 11980 5704 12032 5710
rect 11980 5646 12032 5652
rect 11520 5364 11572 5370
rect 11520 5306 11572 5312
rect 11428 5160 11480 5166
rect 11428 5102 11480 5108
rect 11440 4758 11468 5102
rect 11504 4924 11812 4933
rect 11504 4922 11510 4924
rect 11566 4922 11590 4924
rect 11646 4922 11670 4924
rect 11726 4922 11750 4924
rect 11806 4922 11812 4924
rect 11566 4870 11568 4922
rect 11748 4870 11750 4922
rect 11504 4868 11510 4870
rect 11566 4868 11590 4870
rect 11646 4868 11670 4870
rect 11726 4868 11750 4870
rect 11806 4868 11812 4870
rect 11504 4859 11812 4868
rect 11520 4820 11572 4826
rect 11520 4762 11572 4768
rect 11428 4752 11480 4758
rect 11532 4729 11560 4762
rect 11428 4694 11480 4700
rect 11518 4720 11574 4729
rect 11518 4655 11574 4664
rect 11520 4616 11572 4622
rect 11520 4558 11572 4564
rect 11532 4282 11560 4558
rect 11992 4298 12020 5646
rect 12084 5250 12112 6854
rect 12162 6800 12218 7200
rect 12530 6800 12586 7200
rect 12898 6800 12954 7200
rect 13266 6800 13322 7200
rect 13634 6800 13690 7200
rect 14002 6800 14058 7200
rect 14370 6800 14426 7200
rect 14738 6800 14794 7200
rect 15106 6800 15162 7200
rect 12176 6746 12204 6800
rect 12256 6792 12308 6798
rect 12176 6740 12256 6746
rect 12176 6734 12308 6740
rect 12176 6718 12296 6734
rect 12348 6180 12400 6186
rect 12348 6122 12400 6128
rect 12256 5908 12308 5914
rect 12256 5850 12308 5856
rect 12268 5574 12296 5850
rect 12256 5568 12308 5574
rect 12256 5510 12308 5516
rect 12360 5370 12388 6122
rect 12544 5794 12572 6800
rect 12912 6662 12940 6800
rect 12900 6656 12952 6662
rect 12900 6598 12952 6604
rect 12624 6316 12676 6322
rect 12624 6258 12676 6264
rect 12452 5766 12572 5794
rect 12348 5364 12400 5370
rect 12348 5306 12400 5312
rect 12084 5222 12296 5250
rect 12268 5166 12296 5222
rect 12164 5160 12216 5166
rect 12164 5102 12216 5108
rect 12256 5160 12308 5166
rect 12256 5102 12308 5108
rect 12072 4752 12124 4758
rect 12072 4694 12124 4700
rect 12084 4486 12112 4694
rect 12176 4622 12204 5102
rect 12256 5024 12308 5030
rect 12256 4966 12308 4972
rect 12348 5024 12400 5030
rect 12348 4966 12400 4972
rect 12268 4622 12296 4966
rect 12164 4616 12216 4622
rect 12164 4558 12216 4564
rect 12256 4616 12308 4622
rect 12256 4558 12308 4564
rect 12072 4480 12124 4486
rect 12072 4422 12124 4428
rect 11520 4276 11572 4282
rect 11992 4270 12296 4298
rect 11520 4218 11572 4224
rect 12164 4140 12216 4146
rect 12164 4082 12216 4088
rect 11888 4004 11940 4010
rect 11888 3946 11940 3952
rect 11504 3836 11812 3845
rect 11504 3834 11510 3836
rect 11566 3834 11590 3836
rect 11646 3834 11670 3836
rect 11726 3834 11750 3836
rect 11806 3834 11812 3836
rect 11566 3782 11568 3834
rect 11748 3782 11750 3834
rect 11504 3780 11510 3782
rect 11566 3780 11590 3782
rect 11646 3780 11670 3782
rect 11726 3780 11750 3782
rect 11806 3780 11812 3782
rect 11504 3771 11812 3780
rect 11796 3732 11848 3738
rect 11796 3674 11848 3680
rect 11808 3058 11836 3674
rect 11900 3602 11928 3946
rect 12176 3942 12204 4082
rect 12268 3942 12296 4270
rect 12164 3936 12216 3942
rect 12164 3878 12216 3884
rect 12256 3936 12308 3942
rect 12256 3878 12308 3884
rect 11888 3596 11940 3602
rect 11888 3538 11940 3544
rect 11980 3596 12032 3602
rect 11980 3538 12032 3544
rect 11992 3194 12020 3538
rect 12176 3466 12204 3878
rect 12164 3460 12216 3466
rect 12164 3402 12216 3408
rect 12256 3460 12308 3466
rect 12256 3402 12308 3408
rect 11980 3188 12032 3194
rect 11980 3130 12032 3136
rect 12268 3058 12296 3402
rect 11336 3052 11388 3058
rect 11336 2994 11388 3000
rect 11796 3052 11848 3058
rect 11796 2994 11848 3000
rect 12256 3052 12308 3058
rect 12256 2994 12308 3000
rect 11244 1896 11296 1902
rect 11244 1838 11296 1844
rect 10600 1352 10652 1358
rect 10600 1294 10652 1300
rect 11348 1306 11376 2994
rect 12256 2848 12308 2854
rect 12256 2790 12308 2796
rect 11504 2748 11812 2757
rect 11504 2746 11510 2748
rect 11566 2746 11590 2748
rect 11646 2746 11670 2748
rect 11726 2746 11750 2748
rect 11806 2746 11812 2748
rect 11566 2694 11568 2746
rect 11748 2694 11750 2746
rect 11504 2692 11510 2694
rect 11566 2692 11590 2694
rect 11646 2692 11670 2694
rect 11726 2692 11750 2694
rect 11806 2692 11812 2694
rect 11504 2683 11812 2692
rect 11428 2508 11480 2514
rect 11428 2450 11480 2456
rect 11440 1766 11468 2450
rect 12070 2408 12126 2417
rect 12070 2343 12126 2352
rect 11520 2304 11572 2310
rect 11520 2246 11572 2252
rect 11532 2106 11560 2246
rect 11520 2100 11572 2106
rect 11520 2042 11572 2048
rect 12084 1766 12112 2343
rect 11428 1760 11480 1766
rect 11428 1702 11480 1708
rect 11888 1760 11940 1766
rect 11888 1702 11940 1708
rect 12072 1760 12124 1766
rect 12072 1702 12124 1708
rect 11504 1660 11812 1669
rect 11504 1658 11510 1660
rect 11566 1658 11590 1660
rect 11646 1658 11670 1660
rect 11726 1658 11750 1660
rect 11806 1658 11812 1660
rect 11566 1606 11568 1658
rect 11748 1606 11750 1658
rect 11504 1604 11510 1606
rect 11566 1604 11590 1606
rect 11646 1604 11670 1606
rect 11726 1604 11750 1606
rect 11806 1604 11812 1606
rect 11504 1595 11812 1604
rect 11900 1562 11928 1702
rect 11888 1556 11940 1562
rect 11888 1498 11940 1504
rect 12268 1494 12296 2790
rect 12256 1488 12308 1494
rect 12256 1430 12308 1436
rect 11428 1352 11480 1358
rect 11348 1300 11428 1306
rect 11348 1294 11480 1300
rect 11348 1278 11468 1294
rect 11348 1018 11376 1278
rect 12360 1018 12388 4966
rect 12452 4298 12480 5766
rect 12532 5704 12584 5710
rect 12532 5646 12584 5652
rect 12544 5370 12572 5646
rect 12636 5642 12664 6258
rect 12808 6112 12860 6118
rect 12808 6054 12860 6060
rect 12992 6112 13044 6118
rect 12992 6054 13044 6060
rect 12716 5772 12768 5778
rect 12716 5714 12768 5720
rect 12624 5636 12676 5642
rect 12624 5578 12676 5584
rect 12532 5364 12584 5370
rect 12532 5306 12584 5312
rect 12636 5234 12664 5578
rect 12624 5228 12676 5234
rect 12624 5170 12676 5176
rect 12728 5114 12756 5714
rect 12636 5086 12756 5114
rect 12636 4690 12664 5086
rect 12716 5024 12768 5030
rect 12716 4966 12768 4972
rect 12624 4684 12676 4690
rect 12624 4626 12676 4632
rect 12452 4270 12664 4298
rect 12532 4140 12584 4146
rect 12532 4082 12584 4088
rect 12544 3670 12572 4082
rect 12532 3664 12584 3670
rect 12532 3606 12584 3612
rect 12440 3052 12492 3058
rect 12440 2994 12492 3000
rect 12452 1970 12480 2994
rect 12532 2984 12584 2990
rect 12636 2961 12664 4270
rect 12728 4146 12756 4966
rect 12820 4486 12848 6054
rect 12900 5636 12952 5642
rect 12900 5578 12952 5584
rect 12912 4690 12940 5578
rect 12900 4684 12952 4690
rect 12900 4626 12952 4632
rect 12808 4480 12860 4486
rect 12808 4422 12860 4428
rect 12716 4140 12768 4146
rect 12716 4082 12768 4088
rect 12808 4140 12860 4146
rect 12808 4082 12860 4088
rect 12820 3346 12848 4082
rect 13004 3738 13032 6054
rect 13084 5024 13136 5030
rect 13084 4966 13136 4972
rect 13096 4622 13124 4966
rect 13176 4684 13228 4690
rect 13176 4626 13228 4632
rect 13084 4616 13136 4622
rect 13084 4558 13136 4564
rect 13084 4480 13136 4486
rect 13084 4422 13136 4428
rect 13096 4146 13124 4422
rect 13084 4140 13136 4146
rect 13084 4082 13136 4088
rect 12992 3732 13044 3738
rect 12992 3674 13044 3680
rect 12820 3318 12940 3346
rect 12912 3194 12940 3318
rect 12900 3188 12952 3194
rect 12900 3130 12952 3136
rect 12716 2984 12768 2990
rect 12532 2926 12584 2932
rect 12622 2952 12678 2961
rect 12544 2514 12572 2926
rect 12716 2926 12768 2932
rect 12622 2887 12678 2896
rect 12728 2854 12756 2926
rect 12716 2848 12768 2854
rect 12716 2790 12768 2796
rect 12728 2650 12756 2790
rect 13004 2650 13032 3674
rect 13096 3670 13124 4082
rect 13188 3942 13216 4626
rect 13176 3936 13228 3942
rect 13176 3878 13228 3884
rect 13084 3664 13136 3670
rect 13084 3606 13136 3612
rect 13174 3632 13230 3641
rect 13174 3567 13176 3576
rect 13228 3567 13230 3576
rect 13176 3538 13228 3544
rect 13188 3482 13216 3538
rect 13096 3454 13216 3482
rect 12716 2644 12768 2650
rect 12716 2586 12768 2592
rect 12992 2644 13044 2650
rect 12992 2586 13044 2592
rect 12728 2530 12756 2586
rect 13096 2530 13124 3454
rect 13176 3392 13228 3398
rect 13176 3334 13228 3340
rect 13188 3126 13216 3334
rect 13176 3120 13228 3126
rect 13176 3062 13228 3068
rect 13280 2666 13308 6800
rect 13648 6644 13676 6800
rect 13648 6616 13768 6644
rect 13355 6556 13663 6565
rect 13355 6554 13361 6556
rect 13417 6554 13441 6556
rect 13497 6554 13521 6556
rect 13577 6554 13601 6556
rect 13657 6554 13663 6556
rect 13417 6502 13419 6554
rect 13599 6502 13601 6554
rect 13355 6500 13361 6502
rect 13417 6500 13441 6502
rect 13497 6500 13521 6502
rect 13577 6500 13601 6502
rect 13657 6500 13663 6502
rect 13355 6491 13663 6500
rect 13544 6316 13596 6322
rect 13544 6258 13596 6264
rect 13556 5778 13584 6258
rect 13544 5772 13596 5778
rect 13544 5714 13596 5720
rect 13740 5658 13768 6616
rect 14016 6254 14044 6800
rect 14280 6384 14332 6390
rect 14280 6326 14332 6332
rect 14004 6248 14056 6254
rect 14004 6190 14056 6196
rect 14188 6180 14240 6186
rect 14188 6122 14240 6128
rect 13820 6112 13872 6118
rect 13820 6054 13872 6060
rect 14096 6112 14148 6118
rect 14096 6054 14148 6060
rect 13832 5846 13860 6054
rect 13820 5840 13872 5846
rect 13820 5782 13872 5788
rect 13912 5772 13964 5778
rect 13912 5714 13964 5720
rect 13740 5630 13860 5658
rect 13728 5568 13780 5574
rect 13728 5510 13780 5516
rect 13355 5468 13663 5477
rect 13355 5466 13361 5468
rect 13417 5466 13441 5468
rect 13497 5466 13521 5468
rect 13577 5466 13601 5468
rect 13657 5466 13663 5468
rect 13417 5414 13419 5466
rect 13599 5414 13601 5466
rect 13355 5412 13361 5414
rect 13417 5412 13441 5414
rect 13497 5412 13521 5414
rect 13577 5412 13601 5414
rect 13657 5412 13663 5414
rect 13355 5403 13663 5412
rect 13740 5166 13768 5510
rect 13728 5160 13780 5166
rect 13728 5102 13780 5108
rect 13832 5012 13860 5630
rect 13924 5166 13952 5714
rect 14004 5704 14056 5710
rect 14004 5646 14056 5652
rect 13912 5160 13964 5166
rect 13912 5102 13964 5108
rect 13740 4984 13860 5012
rect 13912 5024 13964 5030
rect 13355 4380 13663 4389
rect 13355 4378 13361 4380
rect 13417 4378 13441 4380
rect 13497 4378 13521 4380
rect 13577 4378 13601 4380
rect 13657 4378 13663 4380
rect 13417 4326 13419 4378
rect 13599 4326 13601 4378
rect 13355 4324 13361 4326
rect 13417 4324 13441 4326
rect 13497 4324 13521 4326
rect 13577 4324 13601 4326
rect 13657 4324 13663 4326
rect 13355 4315 13663 4324
rect 13360 4004 13412 4010
rect 13360 3946 13412 3952
rect 13372 3398 13400 3946
rect 13360 3392 13412 3398
rect 13360 3334 13412 3340
rect 13355 3292 13663 3301
rect 13355 3290 13361 3292
rect 13417 3290 13441 3292
rect 13497 3290 13521 3292
rect 13577 3290 13601 3292
rect 13657 3290 13663 3292
rect 13417 3238 13419 3290
rect 13599 3238 13601 3290
rect 13355 3236 13361 3238
rect 13417 3236 13441 3238
rect 13497 3236 13521 3238
rect 13577 3236 13601 3238
rect 13657 3236 13663 3238
rect 13355 3227 13663 3236
rect 12532 2508 12584 2514
rect 12728 2502 12940 2530
rect 13004 2514 13124 2530
rect 12532 2450 12584 2456
rect 12912 2378 12940 2502
rect 12992 2508 13124 2514
rect 13044 2502 13124 2508
rect 13188 2638 13308 2666
rect 12992 2450 13044 2456
rect 13084 2440 13136 2446
rect 13084 2382 13136 2388
rect 12900 2372 12952 2378
rect 12900 2314 12952 2320
rect 12808 2100 12860 2106
rect 12808 2042 12860 2048
rect 12440 1964 12492 1970
rect 12440 1906 12492 1912
rect 12440 1828 12492 1834
rect 12440 1770 12492 1776
rect 12716 1828 12768 1834
rect 12716 1770 12768 1776
rect 12452 1018 12480 1770
rect 12728 1562 12756 1770
rect 12820 1562 12848 2042
rect 13096 2038 13124 2382
rect 13188 2106 13216 2638
rect 13268 2508 13320 2514
rect 13268 2450 13320 2456
rect 13176 2100 13228 2106
rect 13176 2042 13228 2048
rect 13084 2032 13136 2038
rect 13084 1974 13136 1980
rect 12992 1828 13044 1834
rect 12992 1770 13044 1776
rect 12716 1556 12768 1562
rect 12716 1498 12768 1504
rect 12808 1556 12860 1562
rect 12808 1498 12860 1504
rect 13004 1494 13032 1770
rect 12992 1488 13044 1494
rect 12992 1430 13044 1436
rect 13096 1358 13124 1974
rect 13280 1562 13308 2450
rect 13355 2204 13663 2213
rect 13355 2202 13361 2204
rect 13417 2202 13441 2204
rect 13497 2202 13521 2204
rect 13577 2202 13601 2204
rect 13657 2202 13663 2204
rect 13417 2150 13419 2202
rect 13599 2150 13601 2202
rect 13355 2148 13361 2150
rect 13417 2148 13441 2150
rect 13497 2148 13521 2150
rect 13577 2148 13601 2150
rect 13657 2148 13663 2150
rect 13355 2139 13663 2148
rect 13360 2032 13412 2038
rect 13358 2000 13360 2009
rect 13636 2032 13688 2038
rect 13412 2000 13414 2009
rect 13636 1974 13688 1980
rect 13358 1935 13414 1944
rect 13268 1556 13320 1562
rect 13268 1498 13320 1504
rect 13648 1442 13676 1974
rect 13740 1562 13768 4984
rect 13912 4966 13964 4972
rect 13924 4593 13952 4966
rect 13910 4584 13966 4593
rect 13910 4519 13966 4528
rect 14016 4078 14044 5646
rect 14108 5234 14136 6054
rect 14096 5228 14148 5234
rect 14096 5170 14148 5176
rect 14200 4826 14228 6122
rect 14188 4820 14240 4826
rect 14188 4762 14240 4768
rect 14292 4706 14320 6326
rect 14200 4678 14320 4706
rect 14384 4690 14412 6800
rect 14648 6316 14700 6322
rect 14648 6258 14700 6264
rect 14556 5704 14608 5710
rect 14556 5646 14608 5652
rect 14372 4684 14424 4690
rect 14096 4140 14148 4146
rect 14096 4082 14148 4088
rect 13912 4072 13964 4078
rect 13912 4014 13964 4020
rect 14004 4072 14056 4078
rect 14004 4014 14056 4020
rect 13924 3738 13952 4014
rect 14108 3777 14136 4082
rect 14094 3768 14150 3777
rect 13912 3732 13964 3738
rect 14094 3703 14150 3712
rect 13912 3674 13964 3680
rect 14096 3596 14148 3602
rect 14016 3556 14096 3584
rect 13820 2848 13872 2854
rect 13820 2790 13872 2796
rect 13832 2446 13860 2790
rect 13820 2440 13872 2446
rect 13820 2382 13872 2388
rect 13728 1556 13780 1562
rect 13728 1498 13780 1504
rect 13648 1414 13768 1442
rect 13084 1352 13136 1358
rect 13176 1352 13228 1358
rect 13084 1294 13136 1300
rect 13174 1320 13176 1329
rect 13228 1320 13230 1329
rect 13174 1255 13230 1264
rect 13355 1116 13663 1125
rect 13355 1114 13361 1116
rect 13417 1114 13441 1116
rect 13497 1114 13521 1116
rect 13577 1114 13601 1116
rect 13657 1114 13663 1116
rect 13417 1062 13419 1114
rect 13599 1062 13601 1114
rect 13355 1060 13361 1062
rect 13417 1060 13441 1062
rect 13497 1060 13521 1062
rect 13577 1060 13601 1062
rect 13657 1060 13663 1062
rect 13355 1051 13663 1060
rect 11336 1012 11388 1018
rect 11336 954 11388 960
rect 12348 1012 12400 1018
rect 12348 954 12400 960
rect 12440 1012 12492 1018
rect 12440 954 12492 960
rect 13740 814 13768 1414
rect 13832 1018 13860 2382
rect 14016 1766 14044 3556
rect 14200 3584 14228 4678
rect 14372 4626 14424 4632
rect 14464 4616 14516 4622
rect 14464 4558 14516 4564
rect 14148 3556 14228 3584
rect 14096 3538 14148 3544
rect 14094 3496 14150 3505
rect 14094 3431 14150 3440
rect 14108 3058 14136 3431
rect 14188 3392 14240 3398
rect 14188 3334 14240 3340
rect 14096 3052 14148 3058
rect 14096 2994 14148 3000
rect 14108 2650 14136 2994
rect 14200 2854 14228 3334
rect 14188 2848 14240 2854
rect 14188 2790 14240 2796
rect 14096 2644 14148 2650
rect 14096 2586 14148 2592
rect 14372 2508 14424 2514
rect 14372 2450 14424 2456
rect 14188 2304 14240 2310
rect 14188 2246 14240 2252
rect 14200 1902 14228 2246
rect 14188 1896 14240 1902
rect 14188 1838 14240 1844
rect 14004 1760 14056 1766
rect 14004 1702 14056 1708
rect 14384 1562 14412 2450
rect 14476 2378 14504 4558
rect 14568 4049 14596 5646
rect 14660 4690 14688 6258
rect 14648 4684 14700 4690
rect 14648 4626 14700 4632
rect 14660 4146 14688 4626
rect 14648 4140 14700 4146
rect 14648 4082 14700 4088
rect 14554 4040 14610 4049
rect 14554 3975 14610 3984
rect 14556 3936 14608 3942
rect 14556 3878 14608 3884
rect 14568 2802 14596 3878
rect 14648 3120 14700 3126
rect 14646 3088 14648 3097
rect 14700 3088 14702 3097
rect 14646 3023 14702 3032
rect 14646 2952 14702 2961
rect 14646 2887 14648 2896
rect 14700 2887 14702 2896
rect 14648 2858 14700 2864
rect 14568 2774 14688 2802
rect 14556 2576 14608 2582
rect 14556 2518 14608 2524
rect 14464 2372 14516 2378
rect 14464 2314 14516 2320
rect 14372 1556 14424 1562
rect 14372 1498 14424 1504
rect 13912 1284 13964 1290
rect 13912 1226 13964 1232
rect 13820 1012 13872 1018
rect 13820 954 13872 960
rect 13924 950 13952 1226
rect 14568 1018 14596 2518
rect 14660 1562 14688 2774
rect 14752 1562 14780 6800
rect 15016 6792 15068 6798
rect 15016 6734 15068 6740
rect 14832 6112 14884 6118
rect 14832 6054 14884 6060
rect 14844 5914 14872 6054
rect 14832 5908 14884 5914
rect 14832 5850 14884 5856
rect 14844 3942 14872 5850
rect 14924 5228 14976 5234
rect 14924 5170 14976 5176
rect 14832 3936 14884 3942
rect 14832 3878 14884 3884
rect 14648 1556 14700 1562
rect 14648 1498 14700 1504
rect 14740 1556 14792 1562
rect 14740 1498 14792 1504
rect 14556 1012 14608 1018
rect 14556 954 14608 960
rect 13912 944 13964 950
rect 13912 886 13964 892
rect 940 808 992 814
rect 860 768 940 796
rect 860 400 888 768
rect 1952 808 2004 814
rect 940 750 992 756
rect 1872 768 1952 796
rect 1872 400 1900 768
rect 1952 750 2004 756
rect 2872 808 2924 814
rect 2872 750 2924 756
rect 3976 808 4028 814
rect 3976 750 4028 756
rect 4988 808 5040 814
rect 4988 750 5040 756
rect 6184 808 6236 814
rect 6184 750 6236 756
rect 7012 808 7064 814
rect 7012 750 7064 756
rect 7380 808 7432 814
rect 7380 750 7432 756
rect 7472 808 7524 814
rect 7472 750 7524 756
rect 8208 808 8260 814
rect 8208 750 8260 756
rect 10048 808 10100 814
rect 10048 750 10100 756
rect 10508 808 10560 814
rect 10508 750 10560 756
rect 11060 808 11112 814
rect 11060 750 11112 756
rect 12072 808 12124 814
rect 12072 750 12124 756
rect 13084 808 13136 814
rect 13084 750 13136 756
rect 13728 808 13780 814
rect 13728 750 13780 756
rect 14004 808 14056 814
rect 14004 750 14056 756
rect 2884 400 2912 750
rect 3988 490 4016 750
rect 4100 572 4408 581
rect 4100 570 4106 572
rect 4162 570 4186 572
rect 4242 570 4266 572
rect 4322 570 4346 572
rect 4402 570 4408 572
rect 4162 518 4164 570
rect 4344 518 4346 570
rect 4100 516 4106 518
rect 4162 516 4186 518
rect 4242 516 4266 518
rect 4322 516 4346 518
rect 4402 516 4408 518
rect 4100 507 4408 516
rect 5000 490 5028 750
rect 3896 462 4016 490
rect 4908 462 5028 490
rect 5920 462 6040 490
rect 3896 400 3924 462
rect 4908 400 4936 462
rect 5920 400 5948 462
rect 846 0 902 400
rect 1858 0 1914 400
rect 2870 0 2926 400
rect 3882 0 3938 400
rect 4894 0 4950 400
rect 5906 0 5962 400
rect 6012 354 6040 462
rect 6196 354 6224 750
rect 7024 490 7052 750
rect 7802 572 8110 581
rect 7802 570 7808 572
rect 7864 570 7888 572
rect 7944 570 7968 572
rect 8024 570 8048 572
rect 8104 570 8110 572
rect 7864 518 7866 570
rect 8046 518 8048 570
rect 7802 516 7808 518
rect 7864 516 7888 518
rect 7944 516 7968 518
rect 8024 516 8048 518
rect 8104 516 8110 518
rect 7802 507 8110 516
rect 6932 462 7052 490
rect 8220 474 8248 750
rect 8944 740 8996 746
rect 8944 682 8996 688
rect 8024 468 8076 474
rect 6932 400 6960 462
rect 7944 428 8024 456
rect 7944 400 7972 428
rect 8024 410 8076 416
rect 8208 468 8260 474
rect 8208 410 8260 416
rect 8956 400 8984 682
rect 10060 490 10088 750
rect 11072 490 11100 750
rect 11504 572 11812 581
rect 11504 570 11510 572
rect 11566 570 11590 572
rect 11646 570 11670 572
rect 11726 570 11750 572
rect 11806 570 11812 572
rect 11566 518 11568 570
rect 11748 518 11750 570
rect 11504 516 11510 518
rect 11566 516 11590 518
rect 11646 516 11670 518
rect 11726 516 11750 518
rect 11806 516 11812 518
rect 11504 507 11812 516
rect 12084 490 12112 750
rect 13096 490 13124 750
rect 9968 462 10088 490
rect 10980 462 11100 490
rect 11992 462 12112 490
rect 13004 462 13124 490
rect 9968 400 9996 462
rect 10980 400 11008 462
rect 11992 400 12020 462
rect 13004 400 13032 462
rect 14016 400 14044 750
rect 14936 746 14964 5170
rect 15028 2038 15056 6734
rect 15120 4078 15148 6800
rect 15660 6724 15712 6730
rect 15660 6666 15712 6672
rect 15568 6656 15620 6662
rect 15568 6598 15620 6604
rect 15206 6012 15514 6021
rect 15206 6010 15212 6012
rect 15268 6010 15292 6012
rect 15348 6010 15372 6012
rect 15428 6010 15452 6012
rect 15508 6010 15514 6012
rect 15268 5958 15270 6010
rect 15450 5958 15452 6010
rect 15206 5956 15212 5958
rect 15268 5956 15292 5958
rect 15348 5956 15372 5958
rect 15428 5956 15452 5958
rect 15508 5956 15514 5958
rect 15206 5947 15514 5956
rect 15206 4924 15514 4933
rect 15206 4922 15212 4924
rect 15268 4922 15292 4924
rect 15348 4922 15372 4924
rect 15428 4922 15452 4924
rect 15508 4922 15514 4924
rect 15268 4870 15270 4922
rect 15450 4870 15452 4922
rect 15206 4868 15212 4870
rect 15268 4868 15292 4870
rect 15348 4868 15372 4870
rect 15428 4868 15452 4870
rect 15508 4868 15514 4870
rect 15206 4859 15514 4868
rect 15108 4072 15160 4078
rect 15108 4014 15160 4020
rect 15108 3936 15160 3942
rect 15108 3878 15160 3884
rect 15016 2032 15068 2038
rect 15016 1974 15068 1980
rect 15016 808 15068 814
rect 15016 750 15068 756
rect 14924 740 14976 746
rect 14924 682 14976 688
rect 15028 400 15056 750
rect 15120 678 15148 3878
rect 15206 3836 15514 3845
rect 15206 3834 15212 3836
rect 15268 3834 15292 3836
rect 15348 3834 15372 3836
rect 15428 3834 15452 3836
rect 15508 3834 15514 3836
rect 15268 3782 15270 3834
rect 15450 3782 15452 3834
rect 15206 3780 15212 3782
rect 15268 3780 15292 3782
rect 15348 3780 15372 3782
rect 15428 3780 15452 3782
rect 15508 3780 15514 3782
rect 15206 3771 15514 3780
rect 15580 3058 15608 6598
rect 15568 3052 15620 3058
rect 15568 2994 15620 3000
rect 15672 2774 15700 6666
rect 15206 2748 15514 2757
rect 15206 2746 15212 2748
rect 15268 2746 15292 2748
rect 15348 2746 15372 2748
rect 15428 2746 15452 2748
rect 15508 2746 15514 2748
rect 15268 2694 15270 2746
rect 15450 2694 15452 2746
rect 15206 2692 15212 2694
rect 15268 2692 15292 2694
rect 15348 2692 15372 2694
rect 15428 2692 15452 2694
rect 15508 2692 15514 2694
rect 15206 2683 15514 2692
rect 15580 2746 15700 2774
rect 15580 2106 15608 2746
rect 15568 2100 15620 2106
rect 15568 2042 15620 2048
rect 15206 1660 15514 1669
rect 15206 1658 15212 1660
rect 15268 1658 15292 1660
rect 15348 1658 15372 1660
rect 15428 1658 15452 1660
rect 15508 1658 15514 1660
rect 15268 1606 15270 1658
rect 15450 1606 15452 1658
rect 15206 1604 15212 1606
rect 15268 1604 15292 1606
rect 15348 1604 15372 1606
rect 15428 1604 15452 1606
rect 15508 1604 15514 1606
rect 15206 1595 15514 1604
rect 15108 672 15160 678
rect 15108 614 15160 620
rect 15206 572 15514 581
rect 15206 570 15212 572
rect 15268 570 15292 572
rect 15348 570 15372 572
rect 15428 570 15452 572
rect 15508 570 15514 572
rect 15268 518 15270 570
rect 15450 518 15452 570
rect 15206 516 15212 518
rect 15268 516 15292 518
rect 15348 516 15372 518
rect 15428 516 15452 518
rect 15508 516 15514 518
rect 15206 507 15514 516
rect 6012 326 6224 354
rect 6918 0 6974 400
rect 7930 0 7986 400
rect 8942 0 8998 400
rect 9954 0 10010 400
rect 10966 0 11022 400
rect 11978 0 12034 400
rect 12990 0 13046 400
rect 14002 0 14058 400
rect 15014 0 15070 400
<< via2 >>
rect 2255 6554 2311 6556
rect 2335 6554 2391 6556
rect 2415 6554 2471 6556
rect 2495 6554 2551 6556
rect 2255 6502 2301 6554
rect 2301 6502 2311 6554
rect 2335 6502 2365 6554
rect 2365 6502 2377 6554
rect 2377 6502 2391 6554
rect 2415 6502 2429 6554
rect 2429 6502 2441 6554
rect 2441 6502 2471 6554
rect 2495 6502 2505 6554
rect 2505 6502 2551 6554
rect 2255 6500 2311 6502
rect 2335 6500 2391 6502
rect 2415 6500 2471 6502
rect 2495 6500 2551 6502
rect 2255 5466 2311 5468
rect 2335 5466 2391 5468
rect 2415 5466 2471 5468
rect 2495 5466 2551 5468
rect 2255 5414 2301 5466
rect 2301 5414 2311 5466
rect 2335 5414 2365 5466
rect 2365 5414 2377 5466
rect 2377 5414 2391 5466
rect 2415 5414 2429 5466
rect 2429 5414 2441 5466
rect 2441 5414 2471 5466
rect 2495 5414 2505 5466
rect 2505 5414 2551 5466
rect 2255 5412 2311 5414
rect 2335 5412 2391 5414
rect 2415 5412 2471 5414
rect 2495 5412 2551 5414
rect 2502 4564 2504 4584
rect 2504 4564 2556 4584
rect 2556 4564 2558 4584
rect 2502 4528 2558 4564
rect 2255 4378 2311 4380
rect 2335 4378 2391 4380
rect 2415 4378 2471 4380
rect 2495 4378 2551 4380
rect 2255 4326 2301 4378
rect 2301 4326 2311 4378
rect 2335 4326 2365 4378
rect 2365 4326 2377 4378
rect 2377 4326 2391 4378
rect 2415 4326 2429 4378
rect 2429 4326 2441 4378
rect 2441 4326 2471 4378
rect 2495 4326 2505 4378
rect 2505 4326 2551 4378
rect 2255 4324 2311 4326
rect 2335 4324 2391 4326
rect 2415 4324 2471 4326
rect 2495 4324 2551 4326
rect 2255 3290 2311 3292
rect 2335 3290 2391 3292
rect 2415 3290 2471 3292
rect 2495 3290 2551 3292
rect 2255 3238 2301 3290
rect 2301 3238 2311 3290
rect 2335 3238 2365 3290
rect 2365 3238 2377 3290
rect 2377 3238 2391 3290
rect 2415 3238 2429 3290
rect 2429 3238 2441 3290
rect 2441 3238 2471 3290
rect 2495 3238 2505 3290
rect 2505 3238 2551 3290
rect 2255 3236 2311 3238
rect 2335 3236 2391 3238
rect 2415 3236 2471 3238
rect 2495 3236 2551 3238
rect 2255 2202 2311 2204
rect 2335 2202 2391 2204
rect 2415 2202 2471 2204
rect 2495 2202 2551 2204
rect 2255 2150 2301 2202
rect 2301 2150 2311 2202
rect 2335 2150 2365 2202
rect 2365 2150 2377 2202
rect 2377 2150 2391 2202
rect 2415 2150 2429 2202
rect 2429 2150 2441 2202
rect 2441 2150 2471 2202
rect 2495 2150 2505 2202
rect 2505 2150 2551 2202
rect 2255 2148 2311 2150
rect 2335 2148 2391 2150
rect 2415 2148 2471 2150
rect 2495 2148 2551 2150
rect 2255 1114 2311 1116
rect 2335 1114 2391 1116
rect 2415 1114 2471 1116
rect 2495 1114 2551 1116
rect 2255 1062 2301 1114
rect 2301 1062 2311 1114
rect 2335 1062 2365 1114
rect 2365 1062 2377 1114
rect 2377 1062 2391 1114
rect 2415 1062 2429 1114
rect 2429 1062 2441 1114
rect 2441 1062 2471 1114
rect 2495 1062 2505 1114
rect 2505 1062 2551 1114
rect 2255 1060 2311 1062
rect 2335 1060 2391 1062
rect 2415 1060 2471 1062
rect 2495 1060 2551 1062
rect 5957 6554 6013 6556
rect 6037 6554 6093 6556
rect 6117 6554 6173 6556
rect 6197 6554 6253 6556
rect 5957 6502 6003 6554
rect 6003 6502 6013 6554
rect 6037 6502 6067 6554
rect 6067 6502 6079 6554
rect 6079 6502 6093 6554
rect 6117 6502 6131 6554
rect 6131 6502 6143 6554
rect 6143 6502 6173 6554
rect 6197 6502 6207 6554
rect 6207 6502 6253 6554
rect 5957 6500 6013 6502
rect 6037 6500 6093 6502
rect 6117 6500 6173 6502
rect 6197 6500 6253 6502
rect 4106 6010 4162 6012
rect 4186 6010 4242 6012
rect 4266 6010 4322 6012
rect 4346 6010 4402 6012
rect 4106 5958 4152 6010
rect 4152 5958 4162 6010
rect 4186 5958 4216 6010
rect 4216 5958 4228 6010
rect 4228 5958 4242 6010
rect 4266 5958 4280 6010
rect 4280 5958 4292 6010
rect 4292 5958 4322 6010
rect 4346 5958 4356 6010
rect 4356 5958 4402 6010
rect 4106 5956 4162 5958
rect 4186 5956 4242 5958
rect 4266 5956 4322 5958
rect 4346 5956 4402 5958
rect 4106 4922 4162 4924
rect 4186 4922 4242 4924
rect 4266 4922 4322 4924
rect 4346 4922 4402 4924
rect 4106 4870 4152 4922
rect 4152 4870 4162 4922
rect 4186 4870 4216 4922
rect 4216 4870 4228 4922
rect 4228 4870 4242 4922
rect 4266 4870 4280 4922
rect 4280 4870 4292 4922
rect 4292 4870 4322 4922
rect 4346 4870 4356 4922
rect 4356 4870 4402 4922
rect 4106 4868 4162 4870
rect 4186 4868 4242 4870
rect 4266 4868 4322 4870
rect 4346 4868 4402 4870
rect 4066 4020 4068 4040
rect 4068 4020 4120 4040
rect 4120 4020 4122 4040
rect 3698 2216 3754 2272
rect 4066 3984 4122 4020
rect 4106 3834 4162 3836
rect 4186 3834 4242 3836
rect 4266 3834 4322 3836
rect 4346 3834 4402 3836
rect 4106 3782 4152 3834
rect 4152 3782 4162 3834
rect 4186 3782 4216 3834
rect 4216 3782 4228 3834
rect 4228 3782 4242 3834
rect 4266 3782 4280 3834
rect 4280 3782 4292 3834
rect 4292 3782 4322 3834
rect 4346 3782 4356 3834
rect 4356 3782 4402 3834
rect 4106 3780 4162 3782
rect 4186 3780 4242 3782
rect 4266 3780 4322 3782
rect 4346 3780 4402 3782
rect 4106 2746 4162 2748
rect 4186 2746 4242 2748
rect 4266 2746 4322 2748
rect 4346 2746 4402 2748
rect 4106 2694 4152 2746
rect 4152 2694 4162 2746
rect 4186 2694 4216 2746
rect 4216 2694 4228 2746
rect 4228 2694 4242 2746
rect 4266 2694 4280 2746
rect 4280 2694 4292 2746
rect 4292 2694 4322 2746
rect 4346 2694 4356 2746
rect 4356 2694 4402 2746
rect 4106 2692 4162 2694
rect 4186 2692 4242 2694
rect 4266 2692 4322 2694
rect 4346 2692 4402 2694
rect 4106 1658 4162 1660
rect 4186 1658 4242 1660
rect 4266 1658 4322 1660
rect 4346 1658 4402 1660
rect 4106 1606 4152 1658
rect 4152 1606 4162 1658
rect 4186 1606 4216 1658
rect 4216 1606 4228 1658
rect 4228 1606 4242 1658
rect 4266 1606 4280 1658
rect 4280 1606 4292 1658
rect 4292 1606 4322 1658
rect 4346 1606 4356 1658
rect 4356 1606 4402 1658
rect 4106 1604 4162 1606
rect 4186 1604 4242 1606
rect 4266 1604 4322 1606
rect 4346 1604 4402 1606
rect 5957 5466 6013 5468
rect 6037 5466 6093 5468
rect 6117 5466 6173 5468
rect 6197 5466 6253 5468
rect 5957 5414 6003 5466
rect 6003 5414 6013 5466
rect 6037 5414 6067 5466
rect 6067 5414 6079 5466
rect 6079 5414 6093 5466
rect 6117 5414 6131 5466
rect 6131 5414 6143 5466
rect 6143 5414 6173 5466
rect 6197 5414 6207 5466
rect 6207 5414 6253 5466
rect 5957 5412 6013 5414
rect 6037 5412 6093 5414
rect 6117 5412 6173 5414
rect 6197 5412 6253 5414
rect 5957 4378 6013 4380
rect 6037 4378 6093 4380
rect 6117 4378 6173 4380
rect 6197 4378 6253 4380
rect 5957 4326 6003 4378
rect 6003 4326 6013 4378
rect 6037 4326 6067 4378
rect 6067 4326 6079 4378
rect 6079 4326 6093 4378
rect 6117 4326 6131 4378
rect 6131 4326 6143 4378
rect 6143 4326 6173 4378
rect 6197 4326 6207 4378
rect 6207 4326 6253 4378
rect 5957 4324 6013 4326
rect 6037 4324 6093 4326
rect 6117 4324 6173 4326
rect 6197 4324 6253 4326
rect 5957 3290 6013 3292
rect 6037 3290 6093 3292
rect 6117 3290 6173 3292
rect 6197 3290 6253 3292
rect 5957 3238 6003 3290
rect 6003 3238 6013 3290
rect 6037 3238 6067 3290
rect 6067 3238 6079 3290
rect 6079 3238 6093 3290
rect 6117 3238 6131 3290
rect 6131 3238 6143 3290
rect 6143 3238 6173 3290
rect 6197 3238 6207 3290
rect 6207 3238 6253 3290
rect 5957 3236 6013 3238
rect 6037 3236 6093 3238
rect 6117 3236 6173 3238
rect 6197 3236 6253 3238
rect 5630 2216 5686 2272
rect 5957 2202 6013 2204
rect 6037 2202 6093 2204
rect 6117 2202 6173 2204
rect 6197 2202 6253 2204
rect 5957 2150 6003 2202
rect 6003 2150 6013 2202
rect 6037 2150 6067 2202
rect 6067 2150 6079 2202
rect 6079 2150 6093 2202
rect 6117 2150 6131 2202
rect 6131 2150 6143 2202
rect 6143 2150 6173 2202
rect 6197 2150 6207 2202
rect 6207 2150 6253 2202
rect 5957 2148 6013 2150
rect 6037 2148 6093 2150
rect 6117 2148 6173 2150
rect 6197 2148 6253 2150
rect 6366 4664 6422 4720
rect 6826 3576 6882 3632
rect 6826 1964 6882 2000
rect 6826 1944 6828 1964
rect 6828 1944 6880 1964
rect 6880 1944 6882 1964
rect 7808 6010 7864 6012
rect 7888 6010 7944 6012
rect 7968 6010 8024 6012
rect 8048 6010 8104 6012
rect 7808 5958 7854 6010
rect 7854 5958 7864 6010
rect 7888 5958 7918 6010
rect 7918 5958 7930 6010
rect 7930 5958 7944 6010
rect 7968 5958 7982 6010
rect 7982 5958 7994 6010
rect 7994 5958 8024 6010
rect 8048 5958 8058 6010
rect 8058 5958 8104 6010
rect 7808 5956 7864 5958
rect 7888 5956 7944 5958
rect 7968 5956 8024 5958
rect 8048 5956 8104 5958
rect 5957 1114 6013 1116
rect 6037 1114 6093 1116
rect 6117 1114 6173 1116
rect 6197 1114 6253 1116
rect 5957 1062 6003 1114
rect 6003 1062 6013 1114
rect 6037 1062 6067 1114
rect 6067 1062 6079 1114
rect 6079 1062 6093 1114
rect 6117 1062 6131 1114
rect 6131 1062 6143 1114
rect 6143 1062 6173 1114
rect 6197 1062 6207 1114
rect 6207 1062 6253 1114
rect 5957 1060 6013 1062
rect 6037 1060 6093 1062
rect 6117 1060 6173 1062
rect 6197 1060 6253 1062
rect 7808 4922 7864 4924
rect 7888 4922 7944 4924
rect 7968 4922 8024 4924
rect 8048 4922 8104 4924
rect 7808 4870 7854 4922
rect 7854 4870 7864 4922
rect 7888 4870 7918 4922
rect 7918 4870 7930 4922
rect 7930 4870 7944 4922
rect 7968 4870 7982 4922
rect 7982 4870 7994 4922
rect 7994 4870 8024 4922
rect 8048 4870 8058 4922
rect 8058 4870 8104 4922
rect 7808 4868 7864 4870
rect 7888 4868 7944 4870
rect 7968 4868 8024 4870
rect 8048 4868 8104 4870
rect 7808 3834 7864 3836
rect 7888 3834 7944 3836
rect 7968 3834 8024 3836
rect 8048 3834 8104 3836
rect 7808 3782 7854 3834
rect 7854 3782 7864 3834
rect 7888 3782 7918 3834
rect 7918 3782 7930 3834
rect 7930 3782 7944 3834
rect 7968 3782 7982 3834
rect 7982 3782 7994 3834
rect 7994 3782 8024 3834
rect 8048 3782 8058 3834
rect 8058 3782 8104 3834
rect 7808 3780 7864 3782
rect 7888 3780 7944 3782
rect 7968 3780 8024 3782
rect 8048 3780 8104 3782
rect 7808 2746 7864 2748
rect 7888 2746 7944 2748
rect 7968 2746 8024 2748
rect 8048 2746 8104 2748
rect 7808 2694 7854 2746
rect 7854 2694 7864 2746
rect 7888 2694 7918 2746
rect 7918 2694 7930 2746
rect 7930 2694 7944 2746
rect 7968 2694 7982 2746
rect 7982 2694 7994 2746
rect 7994 2694 8024 2746
rect 8048 2694 8058 2746
rect 8058 2694 8104 2746
rect 7808 2692 7864 2694
rect 7888 2692 7944 2694
rect 7968 2692 8024 2694
rect 8048 2692 8104 2694
rect 8758 4140 8814 4176
rect 8758 4120 8760 4140
rect 8760 4120 8812 4140
rect 8812 4120 8814 4140
rect 8758 3032 8814 3088
rect 9659 6554 9715 6556
rect 9739 6554 9795 6556
rect 9819 6554 9875 6556
rect 9899 6554 9955 6556
rect 9659 6502 9705 6554
rect 9705 6502 9715 6554
rect 9739 6502 9769 6554
rect 9769 6502 9781 6554
rect 9781 6502 9795 6554
rect 9819 6502 9833 6554
rect 9833 6502 9845 6554
rect 9845 6502 9875 6554
rect 9899 6502 9909 6554
rect 9909 6502 9955 6554
rect 9659 6500 9715 6502
rect 9739 6500 9795 6502
rect 9819 6500 9875 6502
rect 9899 6500 9955 6502
rect 9659 5466 9715 5468
rect 9739 5466 9795 5468
rect 9819 5466 9875 5468
rect 9899 5466 9955 5468
rect 9659 5414 9705 5466
rect 9705 5414 9715 5466
rect 9739 5414 9769 5466
rect 9769 5414 9781 5466
rect 9781 5414 9795 5466
rect 9819 5414 9833 5466
rect 9833 5414 9845 5466
rect 9845 5414 9875 5466
rect 9899 5414 9909 5466
rect 9909 5414 9955 5466
rect 9659 5412 9715 5414
rect 9739 5412 9795 5414
rect 9819 5412 9875 5414
rect 9899 5412 9955 5414
rect 10046 4664 10102 4720
rect 9659 4378 9715 4380
rect 9739 4378 9795 4380
rect 9819 4378 9875 4380
rect 9899 4378 9955 4380
rect 9659 4326 9705 4378
rect 9705 4326 9715 4378
rect 9739 4326 9769 4378
rect 9769 4326 9781 4378
rect 9781 4326 9795 4378
rect 9819 4326 9833 4378
rect 9833 4326 9845 4378
rect 9845 4326 9875 4378
rect 9899 4326 9909 4378
rect 9909 4326 9955 4378
rect 9659 4324 9715 4326
rect 9739 4324 9795 4326
rect 9819 4324 9875 4326
rect 9899 4324 9955 4326
rect 9402 4120 9458 4176
rect 9218 3984 9274 4040
rect 8666 2352 8722 2408
rect 9678 3440 9734 3496
rect 9659 3290 9715 3292
rect 9739 3290 9795 3292
rect 9819 3290 9875 3292
rect 9899 3290 9955 3292
rect 9659 3238 9705 3290
rect 9705 3238 9715 3290
rect 9739 3238 9769 3290
rect 9769 3238 9781 3290
rect 9781 3238 9795 3290
rect 9819 3238 9833 3290
rect 9833 3238 9845 3290
rect 9845 3238 9875 3290
rect 9899 3238 9909 3290
rect 9909 3238 9955 3290
rect 9659 3236 9715 3238
rect 9739 3236 9795 3238
rect 9819 3236 9875 3238
rect 9899 3236 9955 3238
rect 9586 3052 9642 3088
rect 9586 3032 9588 3052
rect 9588 3032 9640 3052
rect 9640 3032 9642 3052
rect 9659 2202 9715 2204
rect 9739 2202 9795 2204
rect 9819 2202 9875 2204
rect 9899 2202 9955 2204
rect 9659 2150 9705 2202
rect 9705 2150 9715 2202
rect 9739 2150 9769 2202
rect 9769 2150 9781 2202
rect 9781 2150 9795 2202
rect 9819 2150 9833 2202
rect 9833 2150 9845 2202
rect 9845 2150 9875 2202
rect 9899 2150 9909 2202
rect 9909 2150 9955 2202
rect 9659 2148 9715 2150
rect 9739 2148 9795 2150
rect 9819 2148 9875 2150
rect 9899 2148 9955 2150
rect 7808 1658 7864 1660
rect 7888 1658 7944 1660
rect 7968 1658 8024 1660
rect 8048 1658 8104 1660
rect 7808 1606 7854 1658
rect 7854 1606 7864 1658
rect 7888 1606 7918 1658
rect 7918 1606 7930 1658
rect 7930 1606 7944 1658
rect 7968 1606 7982 1658
rect 7982 1606 7994 1658
rect 7994 1606 8024 1658
rect 8048 1606 8058 1658
rect 8058 1606 8104 1658
rect 7808 1604 7864 1606
rect 7888 1604 7944 1606
rect 7968 1604 8024 1606
rect 8048 1604 8104 1606
rect 9659 1114 9715 1116
rect 9739 1114 9795 1116
rect 9819 1114 9875 1116
rect 9899 1114 9955 1116
rect 9659 1062 9705 1114
rect 9705 1062 9715 1114
rect 9739 1062 9769 1114
rect 9769 1062 9781 1114
rect 9781 1062 9795 1114
rect 9819 1062 9833 1114
rect 9833 1062 9845 1114
rect 9845 1062 9875 1114
rect 9899 1062 9909 1114
rect 9909 1062 9955 1114
rect 9659 1060 9715 1062
rect 9739 1060 9795 1062
rect 9819 1060 9875 1062
rect 9899 1060 9955 1062
rect 10414 3440 10470 3496
rect 11510 6010 11566 6012
rect 11590 6010 11646 6012
rect 11670 6010 11726 6012
rect 11750 6010 11806 6012
rect 11510 5958 11556 6010
rect 11556 5958 11566 6010
rect 11590 5958 11620 6010
rect 11620 5958 11632 6010
rect 11632 5958 11646 6010
rect 11670 5958 11684 6010
rect 11684 5958 11696 6010
rect 11696 5958 11726 6010
rect 11750 5958 11760 6010
rect 11760 5958 11806 6010
rect 11510 5956 11566 5958
rect 11590 5956 11646 5958
rect 11670 5956 11726 5958
rect 11750 5956 11806 5958
rect 10506 3032 10562 3088
rect 11242 3848 11298 3904
rect 11510 4922 11566 4924
rect 11590 4922 11646 4924
rect 11670 4922 11726 4924
rect 11750 4922 11806 4924
rect 11510 4870 11556 4922
rect 11556 4870 11566 4922
rect 11590 4870 11620 4922
rect 11620 4870 11632 4922
rect 11632 4870 11646 4922
rect 11670 4870 11684 4922
rect 11684 4870 11696 4922
rect 11696 4870 11726 4922
rect 11750 4870 11760 4922
rect 11760 4870 11806 4922
rect 11510 4868 11566 4870
rect 11590 4868 11646 4870
rect 11670 4868 11726 4870
rect 11750 4868 11806 4870
rect 11518 4664 11574 4720
rect 11510 3834 11566 3836
rect 11590 3834 11646 3836
rect 11670 3834 11726 3836
rect 11750 3834 11806 3836
rect 11510 3782 11556 3834
rect 11556 3782 11566 3834
rect 11590 3782 11620 3834
rect 11620 3782 11632 3834
rect 11632 3782 11646 3834
rect 11670 3782 11684 3834
rect 11684 3782 11696 3834
rect 11696 3782 11726 3834
rect 11750 3782 11760 3834
rect 11760 3782 11806 3834
rect 11510 3780 11566 3782
rect 11590 3780 11646 3782
rect 11670 3780 11726 3782
rect 11750 3780 11806 3782
rect 11510 2746 11566 2748
rect 11590 2746 11646 2748
rect 11670 2746 11726 2748
rect 11750 2746 11806 2748
rect 11510 2694 11556 2746
rect 11556 2694 11566 2746
rect 11590 2694 11620 2746
rect 11620 2694 11632 2746
rect 11632 2694 11646 2746
rect 11670 2694 11684 2746
rect 11684 2694 11696 2746
rect 11696 2694 11726 2746
rect 11750 2694 11760 2746
rect 11760 2694 11806 2746
rect 11510 2692 11566 2694
rect 11590 2692 11646 2694
rect 11670 2692 11726 2694
rect 11750 2692 11806 2694
rect 12070 2352 12126 2408
rect 11510 1658 11566 1660
rect 11590 1658 11646 1660
rect 11670 1658 11726 1660
rect 11750 1658 11806 1660
rect 11510 1606 11556 1658
rect 11556 1606 11566 1658
rect 11590 1606 11620 1658
rect 11620 1606 11632 1658
rect 11632 1606 11646 1658
rect 11670 1606 11684 1658
rect 11684 1606 11696 1658
rect 11696 1606 11726 1658
rect 11750 1606 11760 1658
rect 11760 1606 11806 1658
rect 11510 1604 11566 1606
rect 11590 1604 11646 1606
rect 11670 1604 11726 1606
rect 11750 1604 11806 1606
rect 12622 2896 12678 2952
rect 13174 3596 13230 3632
rect 13174 3576 13176 3596
rect 13176 3576 13228 3596
rect 13228 3576 13230 3596
rect 13361 6554 13417 6556
rect 13441 6554 13497 6556
rect 13521 6554 13577 6556
rect 13601 6554 13657 6556
rect 13361 6502 13407 6554
rect 13407 6502 13417 6554
rect 13441 6502 13471 6554
rect 13471 6502 13483 6554
rect 13483 6502 13497 6554
rect 13521 6502 13535 6554
rect 13535 6502 13547 6554
rect 13547 6502 13577 6554
rect 13601 6502 13611 6554
rect 13611 6502 13657 6554
rect 13361 6500 13417 6502
rect 13441 6500 13497 6502
rect 13521 6500 13577 6502
rect 13601 6500 13657 6502
rect 13361 5466 13417 5468
rect 13441 5466 13497 5468
rect 13521 5466 13577 5468
rect 13601 5466 13657 5468
rect 13361 5414 13407 5466
rect 13407 5414 13417 5466
rect 13441 5414 13471 5466
rect 13471 5414 13483 5466
rect 13483 5414 13497 5466
rect 13521 5414 13535 5466
rect 13535 5414 13547 5466
rect 13547 5414 13577 5466
rect 13601 5414 13611 5466
rect 13611 5414 13657 5466
rect 13361 5412 13417 5414
rect 13441 5412 13497 5414
rect 13521 5412 13577 5414
rect 13601 5412 13657 5414
rect 13361 4378 13417 4380
rect 13441 4378 13497 4380
rect 13521 4378 13577 4380
rect 13601 4378 13657 4380
rect 13361 4326 13407 4378
rect 13407 4326 13417 4378
rect 13441 4326 13471 4378
rect 13471 4326 13483 4378
rect 13483 4326 13497 4378
rect 13521 4326 13535 4378
rect 13535 4326 13547 4378
rect 13547 4326 13577 4378
rect 13601 4326 13611 4378
rect 13611 4326 13657 4378
rect 13361 4324 13417 4326
rect 13441 4324 13497 4326
rect 13521 4324 13577 4326
rect 13601 4324 13657 4326
rect 13361 3290 13417 3292
rect 13441 3290 13497 3292
rect 13521 3290 13577 3292
rect 13601 3290 13657 3292
rect 13361 3238 13407 3290
rect 13407 3238 13417 3290
rect 13441 3238 13471 3290
rect 13471 3238 13483 3290
rect 13483 3238 13497 3290
rect 13521 3238 13535 3290
rect 13535 3238 13547 3290
rect 13547 3238 13577 3290
rect 13601 3238 13611 3290
rect 13611 3238 13657 3290
rect 13361 3236 13417 3238
rect 13441 3236 13497 3238
rect 13521 3236 13577 3238
rect 13601 3236 13657 3238
rect 13361 2202 13417 2204
rect 13441 2202 13497 2204
rect 13521 2202 13577 2204
rect 13601 2202 13657 2204
rect 13361 2150 13407 2202
rect 13407 2150 13417 2202
rect 13441 2150 13471 2202
rect 13471 2150 13483 2202
rect 13483 2150 13497 2202
rect 13521 2150 13535 2202
rect 13535 2150 13547 2202
rect 13547 2150 13577 2202
rect 13601 2150 13611 2202
rect 13611 2150 13657 2202
rect 13361 2148 13417 2150
rect 13441 2148 13497 2150
rect 13521 2148 13577 2150
rect 13601 2148 13657 2150
rect 13358 1980 13360 2000
rect 13360 1980 13412 2000
rect 13412 1980 13414 2000
rect 13358 1944 13414 1980
rect 13910 4528 13966 4584
rect 14094 3712 14150 3768
rect 13174 1300 13176 1320
rect 13176 1300 13228 1320
rect 13228 1300 13230 1320
rect 13174 1264 13230 1300
rect 13361 1114 13417 1116
rect 13441 1114 13497 1116
rect 13521 1114 13577 1116
rect 13601 1114 13657 1116
rect 13361 1062 13407 1114
rect 13407 1062 13417 1114
rect 13441 1062 13471 1114
rect 13471 1062 13483 1114
rect 13483 1062 13497 1114
rect 13521 1062 13535 1114
rect 13535 1062 13547 1114
rect 13547 1062 13577 1114
rect 13601 1062 13611 1114
rect 13611 1062 13657 1114
rect 13361 1060 13417 1062
rect 13441 1060 13497 1062
rect 13521 1060 13577 1062
rect 13601 1060 13657 1062
rect 14094 3440 14150 3496
rect 14554 3984 14610 4040
rect 14646 3068 14648 3088
rect 14648 3068 14700 3088
rect 14700 3068 14702 3088
rect 14646 3032 14702 3068
rect 14646 2916 14702 2952
rect 14646 2896 14648 2916
rect 14648 2896 14700 2916
rect 14700 2896 14702 2916
rect 4106 570 4162 572
rect 4186 570 4242 572
rect 4266 570 4322 572
rect 4346 570 4402 572
rect 4106 518 4152 570
rect 4152 518 4162 570
rect 4186 518 4216 570
rect 4216 518 4228 570
rect 4228 518 4242 570
rect 4266 518 4280 570
rect 4280 518 4292 570
rect 4292 518 4322 570
rect 4346 518 4356 570
rect 4356 518 4402 570
rect 4106 516 4162 518
rect 4186 516 4242 518
rect 4266 516 4322 518
rect 4346 516 4402 518
rect 7808 570 7864 572
rect 7888 570 7944 572
rect 7968 570 8024 572
rect 8048 570 8104 572
rect 7808 518 7854 570
rect 7854 518 7864 570
rect 7888 518 7918 570
rect 7918 518 7930 570
rect 7930 518 7944 570
rect 7968 518 7982 570
rect 7982 518 7994 570
rect 7994 518 8024 570
rect 8048 518 8058 570
rect 8058 518 8104 570
rect 7808 516 7864 518
rect 7888 516 7944 518
rect 7968 516 8024 518
rect 8048 516 8104 518
rect 11510 570 11566 572
rect 11590 570 11646 572
rect 11670 570 11726 572
rect 11750 570 11806 572
rect 11510 518 11556 570
rect 11556 518 11566 570
rect 11590 518 11620 570
rect 11620 518 11632 570
rect 11632 518 11646 570
rect 11670 518 11684 570
rect 11684 518 11696 570
rect 11696 518 11726 570
rect 11750 518 11760 570
rect 11760 518 11806 570
rect 11510 516 11566 518
rect 11590 516 11646 518
rect 11670 516 11726 518
rect 11750 516 11806 518
rect 15212 6010 15268 6012
rect 15292 6010 15348 6012
rect 15372 6010 15428 6012
rect 15452 6010 15508 6012
rect 15212 5958 15258 6010
rect 15258 5958 15268 6010
rect 15292 5958 15322 6010
rect 15322 5958 15334 6010
rect 15334 5958 15348 6010
rect 15372 5958 15386 6010
rect 15386 5958 15398 6010
rect 15398 5958 15428 6010
rect 15452 5958 15462 6010
rect 15462 5958 15508 6010
rect 15212 5956 15268 5958
rect 15292 5956 15348 5958
rect 15372 5956 15428 5958
rect 15452 5956 15508 5958
rect 15212 4922 15268 4924
rect 15292 4922 15348 4924
rect 15372 4922 15428 4924
rect 15452 4922 15508 4924
rect 15212 4870 15258 4922
rect 15258 4870 15268 4922
rect 15292 4870 15322 4922
rect 15322 4870 15334 4922
rect 15334 4870 15348 4922
rect 15372 4870 15386 4922
rect 15386 4870 15398 4922
rect 15398 4870 15428 4922
rect 15452 4870 15462 4922
rect 15462 4870 15508 4922
rect 15212 4868 15268 4870
rect 15292 4868 15348 4870
rect 15372 4868 15428 4870
rect 15452 4868 15508 4870
rect 15212 3834 15268 3836
rect 15292 3834 15348 3836
rect 15372 3834 15428 3836
rect 15452 3834 15508 3836
rect 15212 3782 15258 3834
rect 15258 3782 15268 3834
rect 15292 3782 15322 3834
rect 15322 3782 15334 3834
rect 15334 3782 15348 3834
rect 15372 3782 15386 3834
rect 15386 3782 15398 3834
rect 15398 3782 15428 3834
rect 15452 3782 15462 3834
rect 15462 3782 15508 3834
rect 15212 3780 15268 3782
rect 15292 3780 15348 3782
rect 15372 3780 15428 3782
rect 15452 3780 15508 3782
rect 15212 2746 15268 2748
rect 15292 2746 15348 2748
rect 15372 2746 15428 2748
rect 15452 2746 15508 2748
rect 15212 2694 15258 2746
rect 15258 2694 15268 2746
rect 15292 2694 15322 2746
rect 15322 2694 15334 2746
rect 15334 2694 15348 2746
rect 15372 2694 15386 2746
rect 15386 2694 15398 2746
rect 15398 2694 15428 2746
rect 15452 2694 15462 2746
rect 15462 2694 15508 2746
rect 15212 2692 15268 2694
rect 15292 2692 15348 2694
rect 15372 2692 15428 2694
rect 15452 2692 15508 2694
rect 15212 1658 15268 1660
rect 15292 1658 15348 1660
rect 15372 1658 15428 1660
rect 15452 1658 15508 1660
rect 15212 1606 15258 1658
rect 15258 1606 15268 1658
rect 15292 1606 15322 1658
rect 15322 1606 15334 1658
rect 15334 1606 15348 1658
rect 15372 1606 15386 1658
rect 15386 1606 15398 1658
rect 15398 1606 15428 1658
rect 15452 1606 15462 1658
rect 15462 1606 15508 1658
rect 15212 1604 15268 1606
rect 15292 1604 15348 1606
rect 15372 1604 15428 1606
rect 15452 1604 15508 1606
rect 15212 570 15268 572
rect 15292 570 15348 572
rect 15372 570 15428 572
rect 15452 570 15508 572
rect 15212 518 15258 570
rect 15258 518 15268 570
rect 15292 518 15322 570
rect 15322 518 15334 570
rect 15334 518 15348 570
rect 15372 518 15386 570
rect 15386 518 15398 570
rect 15398 518 15428 570
rect 15452 518 15462 570
rect 15462 518 15508 570
rect 15212 516 15268 518
rect 15292 516 15348 518
rect 15372 516 15428 518
rect 15452 516 15508 518
<< metal3 >>
rect 2245 6560 2561 6561
rect 2245 6496 2251 6560
rect 2315 6496 2331 6560
rect 2395 6496 2411 6560
rect 2475 6496 2491 6560
rect 2555 6496 2561 6560
rect 2245 6495 2561 6496
rect 5947 6560 6263 6561
rect 5947 6496 5953 6560
rect 6017 6496 6033 6560
rect 6097 6496 6113 6560
rect 6177 6496 6193 6560
rect 6257 6496 6263 6560
rect 5947 6495 6263 6496
rect 9649 6560 9965 6561
rect 9649 6496 9655 6560
rect 9719 6496 9735 6560
rect 9799 6496 9815 6560
rect 9879 6496 9895 6560
rect 9959 6496 9965 6560
rect 9649 6495 9965 6496
rect 13351 6560 13667 6561
rect 13351 6496 13357 6560
rect 13421 6496 13437 6560
rect 13501 6496 13517 6560
rect 13581 6496 13597 6560
rect 13661 6496 13667 6560
rect 13351 6495 13667 6496
rect 4096 6016 4412 6017
rect 4096 5952 4102 6016
rect 4166 5952 4182 6016
rect 4246 5952 4262 6016
rect 4326 5952 4342 6016
rect 4406 5952 4412 6016
rect 4096 5951 4412 5952
rect 7798 6016 8114 6017
rect 7798 5952 7804 6016
rect 7868 5952 7884 6016
rect 7948 5952 7964 6016
rect 8028 5952 8044 6016
rect 8108 5952 8114 6016
rect 7798 5951 8114 5952
rect 11500 6016 11816 6017
rect 11500 5952 11506 6016
rect 11570 5952 11586 6016
rect 11650 5952 11666 6016
rect 11730 5952 11746 6016
rect 11810 5952 11816 6016
rect 11500 5951 11816 5952
rect 15202 6016 15518 6017
rect 15202 5952 15208 6016
rect 15272 5952 15288 6016
rect 15352 5952 15368 6016
rect 15432 5952 15448 6016
rect 15512 5952 15518 6016
rect 15202 5951 15518 5952
rect 2245 5472 2561 5473
rect 2245 5408 2251 5472
rect 2315 5408 2331 5472
rect 2395 5408 2411 5472
rect 2475 5408 2491 5472
rect 2555 5408 2561 5472
rect 2245 5407 2561 5408
rect 5947 5472 6263 5473
rect 5947 5408 5953 5472
rect 6017 5408 6033 5472
rect 6097 5408 6113 5472
rect 6177 5408 6193 5472
rect 6257 5408 6263 5472
rect 5947 5407 6263 5408
rect 9649 5472 9965 5473
rect 9649 5408 9655 5472
rect 9719 5408 9735 5472
rect 9799 5408 9815 5472
rect 9879 5408 9895 5472
rect 9959 5408 9965 5472
rect 9649 5407 9965 5408
rect 13351 5472 13667 5473
rect 13351 5408 13357 5472
rect 13421 5408 13437 5472
rect 13501 5408 13517 5472
rect 13581 5408 13597 5472
rect 13661 5408 13667 5472
rect 13351 5407 13667 5408
rect 4096 4928 4412 4929
rect 4096 4864 4102 4928
rect 4166 4864 4182 4928
rect 4246 4864 4262 4928
rect 4326 4864 4342 4928
rect 4406 4864 4412 4928
rect 4096 4863 4412 4864
rect 7798 4928 8114 4929
rect 7798 4864 7804 4928
rect 7868 4864 7884 4928
rect 7948 4864 7964 4928
rect 8028 4864 8044 4928
rect 8108 4864 8114 4928
rect 7798 4863 8114 4864
rect 11500 4928 11816 4929
rect 11500 4864 11506 4928
rect 11570 4864 11586 4928
rect 11650 4864 11666 4928
rect 11730 4864 11746 4928
rect 11810 4864 11816 4928
rect 11500 4863 11816 4864
rect 15202 4928 15518 4929
rect 15202 4864 15208 4928
rect 15272 4864 15288 4928
rect 15352 4864 15368 4928
rect 15432 4864 15448 4928
rect 15512 4864 15518 4928
rect 15202 4863 15518 4864
rect 6361 4722 6427 4725
rect 10041 4722 10107 4725
rect 11513 4722 11579 4725
rect 6361 4720 11579 4722
rect 6361 4664 6366 4720
rect 6422 4664 10046 4720
rect 10102 4664 11518 4720
rect 11574 4664 11579 4720
rect 6361 4662 11579 4664
rect 6361 4659 6427 4662
rect 10041 4659 10107 4662
rect 11513 4659 11579 4662
rect 2497 4586 2563 4589
rect 13118 4586 13124 4588
rect 2497 4584 13124 4586
rect 2497 4528 2502 4584
rect 2558 4528 13124 4584
rect 2497 4526 13124 4528
rect 2497 4523 2563 4526
rect 13118 4524 13124 4526
rect 13188 4586 13194 4588
rect 13905 4586 13971 4589
rect 13188 4584 13971 4586
rect 13188 4528 13910 4584
rect 13966 4528 13971 4584
rect 13188 4526 13971 4528
rect 13188 4524 13194 4526
rect 13905 4523 13971 4526
rect 2245 4384 2561 4385
rect 2245 4320 2251 4384
rect 2315 4320 2331 4384
rect 2395 4320 2411 4384
rect 2475 4320 2491 4384
rect 2555 4320 2561 4384
rect 2245 4319 2561 4320
rect 5947 4384 6263 4385
rect 5947 4320 5953 4384
rect 6017 4320 6033 4384
rect 6097 4320 6113 4384
rect 6177 4320 6193 4384
rect 6257 4320 6263 4384
rect 5947 4319 6263 4320
rect 9649 4384 9965 4385
rect 9649 4320 9655 4384
rect 9719 4320 9735 4384
rect 9799 4320 9815 4384
rect 9879 4320 9895 4384
rect 9959 4320 9965 4384
rect 9649 4319 9965 4320
rect 13351 4384 13667 4385
rect 13351 4320 13357 4384
rect 13421 4320 13437 4384
rect 13501 4320 13517 4384
rect 13581 4320 13597 4384
rect 13661 4320 13667 4384
rect 13351 4319 13667 4320
rect 8753 4178 8819 4181
rect 9397 4178 9463 4181
rect 8753 4176 9463 4178
rect 8753 4120 8758 4176
rect 8814 4120 9402 4176
rect 9458 4120 9463 4176
rect 8753 4118 9463 4120
rect 8753 4115 8819 4118
rect 9397 4115 9463 4118
rect 4061 4042 4127 4045
rect 9213 4042 9279 4045
rect 14549 4042 14615 4045
rect 4061 4040 9138 4042
rect 4061 3984 4066 4040
rect 4122 3984 9138 4040
rect 4061 3982 9138 3984
rect 4061 3979 4127 3982
rect 9078 3906 9138 3982
rect 9213 4040 14615 4042
rect 9213 3984 9218 4040
rect 9274 3984 14554 4040
rect 14610 3984 14615 4040
rect 9213 3982 14615 3984
rect 9213 3979 9279 3982
rect 14549 3979 14615 3982
rect 11237 3906 11303 3909
rect 9078 3904 11303 3906
rect 9078 3848 11242 3904
rect 11298 3848 11303 3904
rect 9078 3846 11303 3848
rect 11237 3843 11303 3846
rect 4096 3840 4412 3841
rect 4096 3776 4102 3840
rect 4166 3776 4182 3840
rect 4246 3776 4262 3840
rect 4326 3776 4342 3840
rect 4406 3776 4412 3840
rect 4096 3775 4412 3776
rect 7798 3840 8114 3841
rect 7798 3776 7804 3840
rect 7868 3776 7884 3840
rect 7948 3776 7964 3840
rect 8028 3776 8044 3840
rect 8108 3776 8114 3840
rect 7798 3775 8114 3776
rect 11500 3840 11816 3841
rect 11500 3776 11506 3840
rect 11570 3776 11586 3840
rect 11650 3776 11666 3840
rect 11730 3776 11746 3840
rect 11810 3776 11816 3840
rect 11500 3775 11816 3776
rect 15202 3840 15518 3841
rect 15202 3776 15208 3840
rect 15272 3776 15288 3840
rect 15352 3776 15368 3840
rect 15432 3776 15448 3840
rect 15512 3776 15518 3840
rect 15202 3775 15518 3776
rect 14089 3770 14155 3773
rect 14046 3768 14155 3770
rect 14046 3712 14094 3768
rect 14150 3712 14155 3768
rect 14046 3707 14155 3712
rect 6821 3634 6887 3637
rect 13169 3634 13235 3637
rect 6821 3632 13235 3634
rect 6821 3576 6826 3632
rect 6882 3576 13174 3632
rect 13230 3576 13235 3632
rect 6821 3574 13235 3576
rect 6821 3571 6887 3574
rect 13169 3571 13235 3574
rect 14046 3501 14106 3707
rect 9673 3498 9739 3501
rect 10409 3498 10475 3501
rect 9673 3496 10475 3498
rect 9673 3440 9678 3496
rect 9734 3440 10414 3496
rect 10470 3440 10475 3496
rect 9673 3438 10475 3440
rect 14046 3496 14155 3501
rect 14046 3440 14094 3496
rect 14150 3440 14155 3496
rect 14046 3438 14155 3440
rect 9673 3435 9739 3438
rect 10409 3435 10475 3438
rect 14089 3435 14155 3438
rect 2245 3296 2561 3297
rect 2245 3232 2251 3296
rect 2315 3232 2331 3296
rect 2395 3232 2411 3296
rect 2475 3232 2491 3296
rect 2555 3232 2561 3296
rect 2245 3231 2561 3232
rect 5947 3296 6263 3297
rect 5947 3232 5953 3296
rect 6017 3232 6033 3296
rect 6097 3232 6113 3296
rect 6177 3232 6193 3296
rect 6257 3232 6263 3296
rect 5947 3231 6263 3232
rect 9649 3296 9965 3297
rect 9649 3232 9655 3296
rect 9719 3232 9735 3296
rect 9799 3232 9815 3296
rect 9879 3232 9895 3296
rect 9959 3232 9965 3296
rect 9649 3231 9965 3232
rect 13351 3296 13667 3297
rect 13351 3232 13357 3296
rect 13421 3232 13437 3296
rect 13501 3232 13517 3296
rect 13581 3232 13597 3296
rect 13661 3232 13667 3296
rect 13351 3231 13667 3232
rect 8753 3090 8819 3093
rect 9581 3090 9647 3093
rect 8753 3088 9647 3090
rect 8753 3032 8758 3088
rect 8814 3032 9586 3088
rect 9642 3032 9647 3088
rect 8753 3030 9647 3032
rect 8753 3027 8819 3030
rect 9581 3027 9647 3030
rect 10501 3090 10567 3093
rect 14641 3090 14707 3093
rect 10501 3088 14707 3090
rect 10501 3032 10506 3088
rect 10562 3032 14646 3088
rect 14702 3032 14707 3088
rect 10501 3030 14707 3032
rect 10501 3027 10567 3030
rect 14641 3027 14707 3030
rect 12617 2954 12683 2957
rect 14641 2954 14707 2957
rect 12617 2952 14707 2954
rect 12617 2896 12622 2952
rect 12678 2896 14646 2952
rect 14702 2896 14707 2952
rect 12617 2894 14707 2896
rect 12617 2891 12683 2894
rect 14641 2891 14707 2894
rect 4096 2752 4412 2753
rect 4096 2688 4102 2752
rect 4166 2688 4182 2752
rect 4246 2688 4262 2752
rect 4326 2688 4342 2752
rect 4406 2688 4412 2752
rect 4096 2687 4412 2688
rect 7798 2752 8114 2753
rect 7798 2688 7804 2752
rect 7868 2688 7884 2752
rect 7948 2688 7964 2752
rect 8028 2688 8044 2752
rect 8108 2688 8114 2752
rect 7798 2687 8114 2688
rect 11500 2752 11816 2753
rect 11500 2688 11506 2752
rect 11570 2688 11586 2752
rect 11650 2688 11666 2752
rect 11730 2688 11746 2752
rect 11810 2688 11816 2752
rect 11500 2687 11816 2688
rect 15202 2752 15518 2753
rect 15202 2688 15208 2752
rect 15272 2688 15288 2752
rect 15352 2688 15368 2752
rect 15432 2688 15448 2752
rect 15512 2688 15518 2752
rect 15202 2687 15518 2688
rect 8661 2410 8727 2413
rect 12065 2410 12131 2413
rect 8661 2408 12131 2410
rect 8661 2352 8666 2408
rect 8722 2352 12070 2408
rect 12126 2352 12131 2408
rect 8661 2350 12131 2352
rect 8661 2347 8727 2350
rect 12065 2347 12131 2350
rect 3693 2274 3759 2277
rect 5625 2274 5691 2277
rect 3693 2272 5691 2274
rect 3693 2216 3698 2272
rect 3754 2216 5630 2272
rect 5686 2216 5691 2272
rect 3693 2214 5691 2216
rect 3693 2211 3759 2214
rect 5625 2211 5691 2214
rect 2245 2208 2561 2209
rect 2245 2144 2251 2208
rect 2315 2144 2331 2208
rect 2395 2144 2411 2208
rect 2475 2144 2491 2208
rect 2555 2144 2561 2208
rect 2245 2143 2561 2144
rect 5947 2208 6263 2209
rect 5947 2144 5953 2208
rect 6017 2144 6033 2208
rect 6097 2144 6113 2208
rect 6177 2144 6193 2208
rect 6257 2144 6263 2208
rect 5947 2143 6263 2144
rect 9649 2208 9965 2209
rect 9649 2144 9655 2208
rect 9719 2144 9735 2208
rect 9799 2144 9815 2208
rect 9879 2144 9895 2208
rect 9959 2144 9965 2208
rect 9649 2143 9965 2144
rect 13351 2208 13667 2209
rect 13351 2144 13357 2208
rect 13421 2144 13437 2208
rect 13501 2144 13517 2208
rect 13581 2144 13597 2208
rect 13661 2144 13667 2208
rect 13351 2143 13667 2144
rect 6821 2002 6887 2005
rect 13353 2002 13419 2005
rect 6821 2000 13419 2002
rect 6821 1944 6826 2000
rect 6882 1944 13358 2000
rect 13414 1944 13419 2000
rect 6821 1942 13419 1944
rect 6821 1939 6887 1942
rect 13353 1939 13419 1942
rect 4096 1664 4412 1665
rect 4096 1600 4102 1664
rect 4166 1600 4182 1664
rect 4246 1600 4262 1664
rect 4326 1600 4342 1664
rect 4406 1600 4412 1664
rect 4096 1599 4412 1600
rect 7798 1664 8114 1665
rect 7798 1600 7804 1664
rect 7868 1600 7884 1664
rect 7948 1600 7964 1664
rect 8028 1600 8044 1664
rect 8108 1600 8114 1664
rect 7798 1599 8114 1600
rect 11500 1664 11816 1665
rect 11500 1600 11506 1664
rect 11570 1600 11586 1664
rect 11650 1600 11666 1664
rect 11730 1600 11746 1664
rect 11810 1600 11816 1664
rect 11500 1599 11816 1600
rect 15202 1664 15518 1665
rect 15202 1600 15208 1664
rect 15272 1600 15288 1664
rect 15352 1600 15368 1664
rect 15432 1600 15448 1664
rect 15512 1600 15518 1664
rect 15202 1599 15518 1600
rect 13169 1324 13235 1325
rect 13118 1260 13124 1324
rect 13188 1322 13235 1324
rect 13188 1320 13280 1322
rect 13230 1264 13280 1320
rect 13188 1262 13280 1264
rect 13188 1260 13235 1262
rect 13169 1259 13235 1260
rect 2245 1120 2561 1121
rect 2245 1056 2251 1120
rect 2315 1056 2331 1120
rect 2395 1056 2411 1120
rect 2475 1056 2491 1120
rect 2555 1056 2561 1120
rect 2245 1055 2561 1056
rect 5947 1120 6263 1121
rect 5947 1056 5953 1120
rect 6017 1056 6033 1120
rect 6097 1056 6113 1120
rect 6177 1056 6193 1120
rect 6257 1056 6263 1120
rect 5947 1055 6263 1056
rect 9649 1120 9965 1121
rect 9649 1056 9655 1120
rect 9719 1056 9735 1120
rect 9799 1056 9815 1120
rect 9879 1056 9895 1120
rect 9959 1056 9965 1120
rect 9649 1055 9965 1056
rect 13351 1120 13667 1121
rect 13351 1056 13357 1120
rect 13421 1056 13437 1120
rect 13501 1056 13517 1120
rect 13581 1056 13597 1120
rect 13661 1056 13667 1120
rect 13351 1055 13667 1056
rect 4096 576 4412 577
rect 4096 512 4102 576
rect 4166 512 4182 576
rect 4246 512 4262 576
rect 4326 512 4342 576
rect 4406 512 4412 576
rect 4096 511 4412 512
rect 7798 576 8114 577
rect 7798 512 7804 576
rect 7868 512 7884 576
rect 7948 512 7964 576
rect 8028 512 8044 576
rect 8108 512 8114 576
rect 7798 511 8114 512
rect 11500 576 11816 577
rect 11500 512 11506 576
rect 11570 512 11586 576
rect 11650 512 11666 576
rect 11730 512 11746 576
rect 11810 512 11816 576
rect 11500 511 11816 512
rect 15202 576 15518 577
rect 15202 512 15208 576
rect 15272 512 15288 576
rect 15352 512 15368 576
rect 15432 512 15448 576
rect 15512 512 15518 576
rect 15202 511 15518 512
<< via3 >>
rect 2251 6556 2315 6560
rect 2251 6500 2255 6556
rect 2255 6500 2311 6556
rect 2311 6500 2315 6556
rect 2251 6496 2315 6500
rect 2331 6556 2395 6560
rect 2331 6500 2335 6556
rect 2335 6500 2391 6556
rect 2391 6500 2395 6556
rect 2331 6496 2395 6500
rect 2411 6556 2475 6560
rect 2411 6500 2415 6556
rect 2415 6500 2471 6556
rect 2471 6500 2475 6556
rect 2411 6496 2475 6500
rect 2491 6556 2555 6560
rect 2491 6500 2495 6556
rect 2495 6500 2551 6556
rect 2551 6500 2555 6556
rect 2491 6496 2555 6500
rect 5953 6556 6017 6560
rect 5953 6500 5957 6556
rect 5957 6500 6013 6556
rect 6013 6500 6017 6556
rect 5953 6496 6017 6500
rect 6033 6556 6097 6560
rect 6033 6500 6037 6556
rect 6037 6500 6093 6556
rect 6093 6500 6097 6556
rect 6033 6496 6097 6500
rect 6113 6556 6177 6560
rect 6113 6500 6117 6556
rect 6117 6500 6173 6556
rect 6173 6500 6177 6556
rect 6113 6496 6177 6500
rect 6193 6556 6257 6560
rect 6193 6500 6197 6556
rect 6197 6500 6253 6556
rect 6253 6500 6257 6556
rect 6193 6496 6257 6500
rect 9655 6556 9719 6560
rect 9655 6500 9659 6556
rect 9659 6500 9715 6556
rect 9715 6500 9719 6556
rect 9655 6496 9719 6500
rect 9735 6556 9799 6560
rect 9735 6500 9739 6556
rect 9739 6500 9795 6556
rect 9795 6500 9799 6556
rect 9735 6496 9799 6500
rect 9815 6556 9879 6560
rect 9815 6500 9819 6556
rect 9819 6500 9875 6556
rect 9875 6500 9879 6556
rect 9815 6496 9879 6500
rect 9895 6556 9959 6560
rect 9895 6500 9899 6556
rect 9899 6500 9955 6556
rect 9955 6500 9959 6556
rect 9895 6496 9959 6500
rect 13357 6556 13421 6560
rect 13357 6500 13361 6556
rect 13361 6500 13417 6556
rect 13417 6500 13421 6556
rect 13357 6496 13421 6500
rect 13437 6556 13501 6560
rect 13437 6500 13441 6556
rect 13441 6500 13497 6556
rect 13497 6500 13501 6556
rect 13437 6496 13501 6500
rect 13517 6556 13581 6560
rect 13517 6500 13521 6556
rect 13521 6500 13577 6556
rect 13577 6500 13581 6556
rect 13517 6496 13581 6500
rect 13597 6556 13661 6560
rect 13597 6500 13601 6556
rect 13601 6500 13657 6556
rect 13657 6500 13661 6556
rect 13597 6496 13661 6500
rect 4102 6012 4166 6016
rect 4102 5956 4106 6012
rect 4106 5956 4162 6012
rect 4162 5956 4166 6012
rect 4102 5952 4166 5956
rect 4182 6012 4246 6016
rect 4182 5956 4186 6012
rect 4186 5956 4242 6012
rect 4242 5956 4246 6012
rect 4182 5952 4246 5956
rect 4262 6012 4326 6016
rect 4262 5956 4266 6012
rect 4266 5956 4322 6012
rect 4322 5956 4326 6012
rect 4262 5952 4326 5956
rect 4342 6012 4406 6016
rect 4342 5956 4346 6012
rect 4346 5956 4402 6012
rect 4402 5956 4406 6012
rect 4342 5952 4406 5956
rect 7804 6012 7868 6016
rect 7804 5956 7808 6012
rect 7808 5956 7864 6012
rect 7864 5956 7868 6012
rect 7804 5952 7868 5956
rect 7884 6012 7948 6016
rect 7884 5956 7888 6012
rect 7888 5956 7944 6012
rect 7944 5956 7948 6012
rect 7884 5952 7948 5956
rect 7964 6012 8028 6016
rect 7964 5956 7968 6012
rect 7968 5956 8024 6012
rect 8024 5956 8028 6012
rect 7964 5952 8028 5956
rect 8044 6012 8108 6016
rect 8044 5956 8048 6012
rect 8048 5956 8104 6012
rect 8104 5956 8108 6012
rect 8044 5952 8108 5956
rect 11506 6012 11570 6016
rect 11506 5956 11510 6012
rect 11510 5956 11566 6012
rect 11566 5956 11570 6012
rect 11506 5952 11570 5956
rect 11586 6012 11650 6016
rect 11586 5956 11590 6012
rect 11590 5956 11646 6012
rect 11646 5956 11650 6012
rect 11586 5952 11650 5956
rect 11666 6012 11730 6016
rect 11666 5956 11670 6012
rect 11670 5956 11726 6012
rect 11726 5956 11730 6012
rect 11666 5952 11730 5956
rect 11746 6012 11810 6016
rect 11746 5956 11750 6012
rect 11750 5956 11806 6012
rect 11806 5956 11810 6012
rect 11746 5952 11810 5956
rect 15208 6012 15272 6016
rect 15208 5956 15212 6012
rect 15212 5956 15268 6012
rect 15268 5956 15272 6012
rect 15208 5952 15272 5956
rect 15288 6012 15352 6016
rect 15288 5956 15292 6012
rect 15292 5956 15348 6012
rect 15348 5956 15352 6012
rect 15288 5952 15352 5956
rect 15368 6012 15432 6016
rect 15368 5956 15372 6012
rect 15372 5956 15428 6012
rect 15428 5956 15432 6012
rect 15368 5952 15432 5956
rect 15448 6012 15512 6016
rect 15448 5956 15452 6012
rect 15452 5956 15508 6012
rect 15508 5956 15512 6012
rect 15448 5952 15512 5956
rect 2251 5468 2315 5472
rect 2251 5412 2255 5468
rect 2255 5412 2311 5468
rect 2311 5412 2315 5468
rect 2251 5408 2315 5412
rect 2331 5468 2395 5472
rect 2331 5412 2335 5468
rect 2335 5412 2391 5468
rect 2391 5412 2395 5468
rect 2331 5408 2395 5412
rect 2411 5468 2475 5472
rect 2411 5412 2415 5468
rect 2415 5412 2471 5468
rect 2471 5412 2475 5468
rect 2411 5408 2475 5412
rect 2491 5468 2555 5472
rect 2491 5412 2495 5468
rect 2495 5412 2551 5468
rect 2551 5412 2555 5468
rect 2491 5408 2555 5412
rect 5953 5468 6017 5472
rect 5953 5412 5957 5468
rect 5957 5412 6013 5468
rect 6013 5412 6017 5468
rect 5953 5408 6017 5412
rect 6033 5468 6097 5472
rect 6033 5412 6037 5468
rect 6037 5412 6093 5468
rect 6093 5412 6097 5468
rect 6033 5408 6097 5412
rect 6113 5468 6177 5472
rect 6113 5412 6117 5468
rect 6117 5412 6173 5468
rect 6173 5412 6177 5468
rect 6113 5408 6177 5412
rect 6193 5468 6257 5472
rect 6193 5412 6197 5468
rect 6197 5412 6253 5468
rect 6253 5412 6257 5468
rect 6193 5408 6257 5412
rect 9655 5468 9719 5472
rect 9655 5412 9659 5468
rect 9659 5412 9715 5468
rect 9715 5412 9719 5468
rect 9655 5408 9719 5412
rect 9735 5468 9799 5472
rect 9735 5412 9739 5468
rect 9739 5412 9795 5468
rect 9795 5412 9799 5468
rect 9735 5408 9799 5412
rect 9815 5468 9879 5472
rect 9815 5412 9819 5468
rect 9819 5412 9875 5468
rect 9875 5412 9879 5468
rect 9815 5408 9879 5412
rect 9895 5468 9959 5472
rect 9895 5412 9899 5468
rect 9899 5412 9955 5468
rect 9955 5412 9959 5468
rect 9895 5408 9959 5412
rect 13357 5468 13421 5472
rect 13357 5412 13361 5468
rect 13361 5412 13417 5468
rect 13417 5412 13421 5468
rect 13357 5408 13421 5412
rect 13437 5468 13501 5472
rect 13437 5412 13441 5468
rect 13441 5412 13497 5468
rect 13497 5412 13501 5468
rect 13437 5408 13501 5412
rect 13517 5468 13581 5472
rect 13517 5412 13521 5468
rect 13521 5412 13577 5468
rect 13577 5412 13581 5468
rect 13517 5408 13581 5412
rect 13597 5468 13661 5472
rect 13597 5412 13601 5468
rect 13601 5412 13657 5468
rect 13657 5412 13661 5468
rect 13597 5408 13661 5412
rect 4102 4924 4166 4928
rect 4102 4868 4106 4924
rect 4106 4868 4162 4924
rect 4162 4868 4166 4924
rect 4102 4864 4166 4868
rect 4182 4924 4246 4928
rect 4182 4868 4186 4924
rect 4186 4868 4242 4924
rect 4242 4868 4246 4924
rect 4182 4864 4246 4868
rect 4262 4924 4326 4928
rect 4262 4868 4266 4924
rect 4266 4868 4322 4924
rect 4322 4868 4326 4924
rect 4262 4864 4326 4868
rect 4342 4924 4406 4928
rect 4342 4868 4346 4924
rect 4346 4868 4402 4924
rect 4402 4868 4406 4924
rect 4342 4864 4406 4868
rect 7804 4924 7868 4928
rect 7804 4868 7808 4924
rect 7808 4868 7864 4924
rect 7864 4868 7868 4924
rect 7804 4864 7868 4868
rect 7884 4924 7948 4928
rect 7884 4868 7888 4924
rect 7888 4868 7944 4924
rect 7944 4868 7948 4924
rect 7884 4864 7948 4868
rect 7964 4924 8028 4928
rect 7964 4868 7968 4924
rect 7968 4868 8024 4924
rect 8024 4868 8028 4924
rect 7964 4864 8028 4868
rect 8044 4924 8108 4928
rect 8044 4868 8048 4924
rect 8048 4868 8104 4924
rect 8104 4868 8108 4924
rect 8044 4864 8108 4868
rect 11506 4924 11570 4928
rect 11506 4868 11510 4924
rect 11510 4868 11566 4924
rect 11566 4868 11570 4924
rect 11506 4864 11570 4868
rect 11586 4924 11650 4928
rect 11586 4868 11590 4924
rect 11590 4868 11646 4924
rect 11646 4868 11650 4924
rect 11586 4864 11650 4868
rect 11666 4924 11730 4928
rect 11666 4868 11670 4924
rect 11670 4868 11726 4924
rect 11726 4868 11730 4924
rect 11666 4864 11730 4868
rect 11746 4924 11810 4928
rect 11746 4868 11750 4924
rect 11750 4868 11806 4924
rect 11806 4868 11810 4924
rect 11746 4864 11810 4868
rect 15208 4924 15272 4928
rect 15208 4868 15212 4924
rect 15212 4868 15268 4924
rect 15268 4868 15272 4924
rect 15208 4864 15272 4868
rect 15288 4924 15352 4928
rect 15288 4868 15292 4924
rect 15292 4868 15348 4924
rect 15348 4868 15352 4924
rect 15288 4864 15352 4868
rect 15368 4924 15432 4928
rect 15368 4868 15372 4924
rect 15372 4868 15428 4924
rect 15428 4868 15432 4924
rect 15368 4864 15432 4868
rect 15448 4924 15512 4928
rect 15448 4868 15452 4924
rect 15452 4868 15508 4924
rect 15508 4868 15512 4924
rect 15448 4864 15512 4868
rect 13124 4524 13188 4588
rect 2251 4380 2315 4384
rect 2251 4324 2255 4380
rect 2255 4324 2311 4380
rect 2311 4324 2315 4380
rect 2251 4320 2315 4324
rect 2331 4380 2395 4384
rect 2331 4324 2335 4380
rect 2335 4324 2391 4380
rect 2391 4324 2395 4380
rect 2331 4320 2395 4324
rect 2411 4380 2475 4384
rect 2411 4324 2415 4380
rect 2415 4324 2471 4380
rect 2471 4324 2475 4380
rect 2411 4320 2475 4324
rect 2491 4380 2555 4384
rect 2491 4324 2495 4380
rect 2495 4324 2551 4380
rect 2551 4324 2555 4380
rect 2491 4320 2555 4324
rect 5953 4380 6017 4384
rect 5953 4324 5957 4380
rect 5957 4324 6013 4380
rect 6013 4324 6017 4380
rect 5953 4320 6017 4324
rect 6033 4380 6097 4384
rect 6033 4324 6037 4380
rect 6037 4324 6093 4380
rect 6093 4324 6097 4380
rect 6033 4320 6097 4324
rect 6113 4380 6177 4384
rect 6113 4324 6117 4380
rect 6117 4324 6173 4380
rect 6173 4324 6177 4380
rect 6113 4320 6177 4324
rect 6193 4380 6257 4384
rect 6193 4324 6197 4380
rect 6197 4324 6253 4380
rect 6253 4324 6257 4380
rect 6193 4320 6257 4324
rect 9655 4380 9719 4384
rect 9655 4324 9659 4380
rect 9659 4324 9715 4380
rect 9715 4324 9719 4380
rect 9655 4320 9719 4324
rect 9735 4380 9799 4384
rect 9735 4324 9739 4380
rect 9739 4324 9795 4380
rect 9795 4324 9799 4380
rect 9735 4320 9799 4324
rect 9815 4380 9879 4384
rect 9815 4324 9819 4380
rect 9819 4324 9875 4380
rect 9875 4324 9879 4380
rect 9815 4320 9879 4324
rect 9895 4380 9959 4384
rect 9895 4324 9899 4380
rect 9899 4324 9955 4380
rect 9955 4324 9959 4380
rect 9895 4320 9959 4324
rect 13357 4380 13421 4384
rect 13357 4324 13361 4380
rect 13361 4324 13417 4380
rect 13417 4324 13421 4380
rect 13357 4320 13421 4324
rect 13437 4380 13501 4384
rect 13437 4324 13441 4380
rect 13441 4324 13497 4380
rect 13497 4324 13501 4380
rect 13437 4320 13501 4324
rect 13517 4380 13581 4384
rect 13517 4324 13521 4380
rect 13521 4324 13577 4380
rect 13577 4324 13581 4380
rect 13517 4320 13581 4324
rect 13597 4380 13661 4384
rect 13597 4324 13601 4380
rect 13601 4324 13657 4380
rect 13657 4324 13661 4380
rect 13597 4320 13661 4324
rect 4102 3836 4166 3840
rect 4102 3780 4106 3836
rect 4106 3780 4162 3836
rect 4162 3780 4166 3836
rect 4102 3776 4166 3780
rect 4182 3836 4246 3840
rect 4182 3780 4186 3836
rect 4186 3780 4242 3836
rect 4242 3780 4246 3836
rect 4182 3776 4246 3780
rect 4262 3836 4326 3840
rect 4262 3780 4266 3836
rect 4266 3780 4322 3836
rect 4322 3780 4326 3836
rect 4262 3776 4326 3780
rect 4342 3836 4406 3840
rect 4342 3780 4346 3836
rect 4346 3780 4402 3836
rect 4402 3780 4406 3836
rect 4342 3776 4406 3780
rect 7804 3836 7868 3840
rect 7804 3780 7808 3836
rect 7808 3780 7864 3836
rect 7864 3780 7868 3836
rect 7804 3776 7868 3780
rect 7884 3836 7948 3840
rect 7884 3780 7888 3836
rect 7888 3780 7944 3836
rect 7944 3780 7948 3836
rect 7884 3776 7948 3780
rect 7964 3836 8028 3840
rect 7964 3780 7968 3836
rect 7968 3780 8024 3836
rect 8024 3780 8028 3836
rect 7964 3776 8028 3780
rect 8044 3836 8108 3840
rect 8044 3780 8048 3836
rect 8048 3780 8104 3836
rect 8104 3780 8108 3836
rect 8044 3776 8108 3780
rect 11506 3836 11570 3840
rect 11506 3780 11510 3836
rect 11510 3780 11566 3836
rect 11566 3780 11570 3836
rect 11506 3776 11570 3780
rect 11586 3836 11650 3840
rect 11586 3780 11590 3836
rect 11590 3780 11646 3836
rect 11646 3780 11650 3836
rect 11586 3776 11650 3780
rect 11666 3836 11730 3840
rect 11666 3780 11670 3836
rect 11670 3780 11726 3836
rect 11726 3780 11730 3836
rect 11666 3776 11730 3780
rect 11746 3836 11810 3840
rect 11746 3780 11750 3836
rect 11750 3780 11806 3836
rect 11806 3780 11810 3836
rect 11746 3776 11810 3780
rect 15208 3836 15272 3840
rect 15208 3780 15212 3836
rect 15212 3780 15268 3836
rect 15268 3780 15272 3836
rect 15208 3776 15272 3780
rect 15288 3836 15352 3840
rect 15288 3780 15292 3836
rect 15292 3780 15348 3836
rect 15348 3780 15352 3836
rect 15288 3776 15352 3780
rect 15368 3836 15432 3840
rect 15368 3780 15372 3836
rect 15372 3780 15428 3836
rect 15428 3780 15432 3836
rect 15368 3776 15432 3780
rect 15448 3836 15512 3840
rect 15448 3780 15452 3836
rect 15452 3780 15508 3836
rect 15508 3780 15512 3836
rect 15448 3776 15512 3780
rect 2251 3292 2315 3296
rect 2251 3236 2255 3292
rect 2255 3236 2311 3292
rect 2311 3236 2315 3292
rect 2251 3232 2315 3236
rect 2331 3292 2395 3296
rect 2331 3236 2335 3292
rect 2335 3236 2391 3292
rect 2391 3236 2395 3292
rect 2331 3232 2395 3236
rect 2411 3292 2475 3296
rect 2411 3236 2415 3292
rect 2415 3236 2471 3292
rect 2471 3236 2475 3292
rect 2411 3232 2475 3236
rect 2491 3292 2555 3296
rect 2491 3236 2495 3292
rect 2495 3236 2551 3292
rect 2551 3236 2555 3292
rect 2491 3232 2555 3236
rect 5953 3292 6017 3296
rect 5953 3236 5957 3292
rect 5957 3236 6013 3292
rect 6013 3236 6017 3292
rect 5953 3232 6017 3236
rect 6033 3292 6097 3296
rect 6033 3236 6037 3292
rect 6037 3236 6093 3292
rect 6093 3236 6097 3292
rect 6033 3232 6097 3236
rect 6113 3292 6177 3296
rect 6113 3236 6117 3292
rect 6117 3236 6173 3292
rect 6173 3236 6177 3292
rect 6113 3232 6177 3236
rect 6193 3292 6257 3296
rect 6193 3236 6197 3292
rect 6197 3236 6253 3292
rect 6253 3236 6257 3292
rect 6193 3232 6257 3236
rect 9655 3292 9719 3296
rect 9655 3236 9659 3292
rect 9659 3236 9715 3292
rect 9715 3236 9719 3292
rect 9655 3232 9719 3236
rect 9735 3292 9799 3296
rect 9735 3236 9739 3292
rect 9739 3236 9795 3292
rect 9795 3236 9799 3292
rect 9735 3232 9799 3236
rect 9815 3292 9879 3296
rect 9815 3236 9819 3292
rect 9819 3236 9875 3292
rect 9875 3236 9879 3292
rect 9815 3232 9879 3236
rect 9895 3292 9959 3296
rect 9895 3236 9899 3292
rect 9899 3236 9955 3292
rect 9955 3236 9959 3292
rect 9895 3232 9959 3236
rect 13357 3292 13421 3296
rect 13357 3236 13361 3292
rect 13361 3236 13417 3292
rect 13417 3236 13421 3292
rect 13357 3232 13421 3236
rect 13437 3292 13501 3296
rect 13437 3236 13441 3292
rect 13441 3236 13497 3292
rect 13497 3236 13501 3292
rect 13437 3232 13501 3236
rect 13517 3292 13581 3296
rect 13517 3236 13521 3292
rect 13521 3236 13577 3292
rect 13577 3236 13581 3292
rect 13517 3232 13581 3236
rect 13597 3292 13661 3296
rect 13597 3236 13601 3292
rect 13601 3236 13657 3292
rect 13657 3236 13661 3292
rect 13597 3232 13661 3236
rect 4102 2748 4166 2752
rect 4102 2692 4106 2748
rect 4106 2692 4162 2748
rect 4162 2692 4166 2748
rect 4102 2688 4166 2692
rect 4182 2748 4246 2752
rect 4182 2692 4186 2748
rect 4186 2692 4242 2748
rect 4242 2692 4246 2748
rect 4182 2688 4246 2692
rect 4262 2748 4326 2752
rect 4262 2692 4266 2748
rect 4266 2692 4322 2748
rect 4322 2692 4326 2748
rect 4262 2688 4326 2692
rect 4342 2748 4406 2752
rect 4342 2692 4346 2748
rect 4346 2692 4402 2748
rect 4402 2692 4406 2748
rect 4342 2688 4406 2692
rect 7804 2748 7868 2752
rect 7804 2692 7808 2748
rect 7808 2692 7864 2748
rect 7864 2692 7868 2748
rect 7804 2688 7868 2692
rect 7884 2748 7948 2752
rect 7884 2692 7888 2748
rect 7888 2692 7944 2748
rect 7944 2692 7948 2748
rect 7884 2688 7948 2692
rect 7964 2748 8028 2752
rect 7964 2692 7968 2748
rect 7968 2692 8024 2748
rect 8024 2692 8028 2748
rect 7964 2688 8028 2692
rect 8044 2748 8108 2752
rect 8044 2692 8048 2748
rect 8048 2692 8104 2748
rect 8104 2692 8108 2748
rect 8044 2688 8108 2692
rect 11506 2748 11570 2752
rect 11506 2692 11510 2748
rect 11510 2692 11566 2748
rect 11566 2692 11570 2748
rect 11506 2688 11570 2692
rect 11586 2748 11650 2752
rect 11586 2692 11590 2748
rect 11590 2692 11646 2748
rect 11646 2692 11650 2748
rect 11586 2688 11650 2692
rect 11666 2748 11730 2752
rect 11666 2692 11670 2748
rect 11670 2692 11726 2748
rect 11726 2692 11730 2748
rect 11666 2688 11730 2692
rect 11746 2748 11810 2752
rect 11746 2692 11750 2748
rect 11750 2692 11806 2748
rect 11806 2692 11810 2748
rect 11746 2688 11810 2692
rect 15208 2748 15272 2752
rect 15208 2692 15212 2748
rect 15212 2692 15268 2748
rect 15268 2692 15272 2748
rect 15208 2688 15272 2692
rect 15288 2748 15352 2752
rect 15288 2692 15292 2748
rect 15292 2692 15348 2748
rect 15348 2692 15352 2748
rect 15288 2688 15352 2692
rect 15368 2748 15432 2752
rect 15368 2692 15372 2748
rect 15372 2692 15428 2748
rect 15428 2692 15432 2748
rect 15368 2688 15432 2692
rect 15448 2748 15512 2752
rect 15448 2692 15452 2748
rect 15452 2692 15508 2748
rect 15508 2692 15512 2748
rect 15448 2688 15512 2692
rect 2251 2204 2315 2208
rect 2251 2148 2255 2204
rect 2255 2148 2311 2204
rect 2311 2148 2315 2204
rect 2251 2144 2315 2148
rect 2331 2204 2395 2208
rect 2331 2148 2335 2204
rect 2335 2148 2391 2204
rect 2391 2148 2395 2204
rect 2331 2144 2395 2148
rect 2411 2204 2475 2208
rect 2411 2148 2415 2204
rect 2415 2148 2471 2204
rect 2471 2148 2475 2204
rect 2411 2144 2475 2148
rect 2491 2204 2555 2208
rect 2491 2148 2495 2204
rect 2495 2148 2551 2204
rect 2551 2148 2555 2204
rect 2491 2144 2555 2148
rect 5953 2204 6017 2208
rect 5953 2148 5957 2204
rect 5957 2148 6013 2204
rect 6013 2148 6017 2204
rect 5953 2144 6017 2148
rect 6033 2204 6097 2208
rect 6033 2148 6037 2204
rect 6037 2148 6093 2204
rect 6093 2148 6097 2204
rect 6033 2144 6097 2148
rect 6113 2204 6177 2208
rect 6113 2148 6117 2204
rect 6117 2148 6173 2204
rect 6173 2148 6177 2204
rect 6113 2144 6177 2148
rect 6193 2204 6257 2208
rect 6193 2148 6197 2204
rect 6197 2148 6253 2204
rect 6253 2148 6257 2204
rect 6193 2144 6257 2148
rect 9655 2204 9719 2208
rect 9655 2148 9659 2204
rect 9659 2148 9715 2204
rect 9715 2148 9719 2204
rect 9655 2144 9719 2148
rect 9735 2204 9799 2208
rect 9735 2148 9739 2204
rect 9739 2148 9795 2204
rect 9795 2148 9799 2204
rect 9735 2144 9799 2148
rect 9815 2204 9879 2208
rect 9815 2148 9819 2204
rect 9819 2148 9875 2204
rect 9875 2148 9879 2204
rect 9815 2144 9879 2148
rect 9895 2204 9959 2208
rect 9895 2148 9899 2204
rect 9899 2148 9955 2204
rect 9955 2148 9959 2204
rect 9895 2144 9959 2148
rect 13357 2204 13421 2208
rect 13357 2148 13361 2204
rect 13361 2148 13417 2204
rect 13417 2148 13421 2204
rect 13357 2144 13421 2148
rect 13437 2204 13501 2208
rect 13437 2148 13441 2204
rect 13441 2148 13497 2204
rect 13497 2148 13501 2204
rect 13437 2144 13501 2148
rect 13517 2204 13581 2208
rect 13517 2148 13521 2204
rect 13521 2148 13577 2204
rect 13577 2148 13581 2204
rect 13517 2144 13581 2148
rect 13597 2204 13661 2208
rect 13597 2148 13601 2204
rect 13601 2148 13657 2204
rect 13657 2148 13661 2204
rect 13597 2144 13661 2148
rect 4102 1660 4166 1664
rect 4102 1604 4106 1660
rect 4106 1604 4162 1660
rect 4162 1604 4166 1660
rect 4102 1600 4166 1604
rect 4182 1660 4246 1664
rect 4182 1604 4186 1660
rect 4186 1604 4242 1660
rect 4242 1604 4246 1660
rect 4182 1600 4246 1604
rect 4262 1660 4326 1664
rect 4262 1604 4266 1660
rect 4266 1604 4322 1660
rect 4322 1604 4326 1660
rect 4262 1600 4326 1604
rect 4342 1660 4406 1664
rect 4342 1604 4346 1660
rect 4346 1604 4402 1660
rect 4402 1604 4406 1660
rect 4342 1600 4406 1604
rect 7804 1660 7868 1664
rect 7804 1604 7808 1660
rect 7808 1604 7864 1660
rect 7864 1604 7868 1660
rect 7804 1600 7868 1604
rect 7884 1660 7948 1664
rect 7884 1604 7888 1660
rect 7888 1604 7944 1660
rect 7944 1604 7948 1660
rect 7884 1600 7948 1604
rect 7964 1660 8028 1664
rect 7964 1604 7968 1660
rect 7968 1604 8024 1660
rect 8024 1604 8028 1660
rect 7964 1600 8028 1604
rect 8044 1660 8108 1664
rect 8044 1604 8048 1660
rect 8048 1604 8104 1660
rect 8104 1604 8108 1660
rect 8044 1600 8108 1604
rect 11506 1660 11570 1664
rect 11506 1604 11510 1660
rect 11510 1604 11566 1660
rect 11566 1604 11570 1660
rect 11506 1600 11570 1604
rect 11586 1660 11650 1664
rect 11586 1604 11590 1660
rect 11590 1604 11646 1660
rect 11646 1604 11650 1660
rect 11586 1600 11650 1604
rect 11666 1660 11730 1664
rect 11666 1604 11670 1660
rect 11670 1604 11726 1660
rect 11726 1604 11730 1660
rect 11666 1600 11730 1604
rect 11746 1660 11810 1664
rect 11746 1604 11750 1660
rect 11750 1604 11806 1660
rect 11806 1604 11810 1660
rect 11746 1600 11810 1604
rect 15208 1660 15272 1664
rect 15208 1604 15212 1660
rect 15212 1604 15268 1660
rect 15268 1604 15272 1660
rect 15208 1600 15272 1604
rect 15288 1660 15352 1664
rect 15288 1604 15292 1660
rect 15292 1604 15348 1660
rect 15348 1604 15352 1660
rect 15288 1600 15352 1604
rect 15368 1660 15432 1664
rect 15368 1604 15372 1660
rect 15372 1604 15428 1660
rect 15428 1604 15432 1660
rect 15368 1600 15432 1604
rect 15448 1660 15512 1664
rect 15448 1604 15452 1660
rect 15452 1604 15508 1660
rect 15508 1604 15512 1660
rect 15448 1600 15512 1604
rect 13124 1320 13188 1324
rect 13124 1264 13174 1320
rect 13174 1264 13188 1320
rect 13124 1260 13188 1264
rect 2251 1116 2315 1120
rect 2251 1060 2255 1116
rect 2255 1060 2311 1116
rect 2311 1060 2315 1116
rect 2251 1056 2315 1060
rect 2331 1116 2395 1120
rect 2331 1060 2335 1116
rect 2335 1060 2391 1116
rect 2391 1060 2395 1116
rect 2331 1056 2395 1060
rect 2411 1116 2475 1120
rect 2411 1060 2415 1116
rect 2415 1060 2471 1116
rect 2471 1060 2475 1116
rect 2411 1056 2475 1060
rect 2491 1116 2555 1120
rect 2491 1060 2495 1116
rect 2495 1060 2551 1116
rect 2551 1060 2555 1116
rect 2491 1056 2555 1060
rect 5953 1116 6017 1120
rect 5953 1060 5957 1116
rect 5957 1060 6013 1116
rect 6013 1060 6017 1116
rect 5953 1056 6017 1060
rect 6033 1116 6097 1120
rect 6033 1060 6037 1116
rect 6037 1060 6093 1116
rect 6093 1060 6097 1116
rect 6033 1056 6097 1060
rect 6113 1116 6177 1120
rect 6113 1060 6117 1116
rect 6117 1060 6173 1116
rect 6173 1060 6177 1116
rect 6113 1056 6177 1060
rect 6193 1116 6257 1120
rect 6193 1060 6197 1116
rect 6197 1060 6253 1116
rect 6253 1060 6257 1116
rect 6193 1056 6257 1060
rect 9655 1116 9719 1120
rect 9655 1060 9659 1116
rect 9659 1060 9715 1116
rect 9715 1060 9719 1116
rect 9655 1056 9719 1060
rect 9735 1116 9799 1120
rect 9735 1060 9739 1116
rect 9739 1060 9795 1116
rect 9795 1060 9799 1116
rect 9735 1056 9799 1060
rect 9815 1116 9879 1120
rect 9815 1060 9819 1116
rect 9819 1060 9875 1116
rect 9875 1060 9879 1116
rect 9815 1056 9879 1060
rect 9895 1116 9959 1120
rect 9895 1060 9899 1116
rect 9899 1060 9955 1116
rect 9955 1060 9959 1116
rect 9895 1056 9959 1060
rect 13357 1116 13421 1120
rect 13357 1060 13361 1116
rect 13361 1060 13417 1116
rect 13417 1060 13421 1116
rect 13357 1056 13421 1060
rect 13437 1116 13501 1120
rect 13437 1060 13441 1116
rect 13441 1060 13497 1116
rect 13497 1060 13501 1116
rect 13437 1056 13501 1060
rect 13517 1116 13581 1120
rect 13517 1060 13521 1116
rect 13521 1060 13577 1116
rect 13577 1060 13581 1116
rect 13517 1056 13581 1060
rect 13597 1116 13661 1120
rect 13597 1060 13601 1116
rect 13601 1060 13657 1116
rect 13657 1060 13661 1116
rect 13597 1056 13661 1060
rect 4102 572 4166 576
rect 4102 516 4106 572
rect 4106 516 4162 572
rect 4162 516 4166 572
rect 4102 512 4166 516
rect 4182 572 4246 576
rect 4182 516 4186 572
rect 4186 516 4242 572
rect 4242 516 4246 572
rect 4182 512 4246 516
rect 4262 572 4326 576
rect 4262 516 4266 572
rect 4266 516 4322 572
rect 4322 516 4326 572
rect 4262 512 4326 516
rect 4342 572 4406 576
rect 4342 516 4346 572
rect 4346 516 4402 572
rect 4402 516 4406 572
rect 4342 512 4406 516
rect 7804 572 7868 576
rect 7804 516 7808 572
rect 7808 516 7864 572
rect 7864 516 7868 572
rect 7804 512 7868 516
rect 7884 572 7948 576
rect 7884 516 7888 572
rect 7888 516 7944 572
rect 7944 516 7948 572
rect 7884 512 7948 516
rect 7964 572 8028 576
rect 7964 516 7968 572
rect 7968 516 8024 572
rect 8024 516 8028 572
rect 7964 512 8028 516
rect 8044 572 8108 576
rect 8044 516 8048 572
rect 8048 516 8104 572
rect 8104 516 8108 572
rect 8044 512 8108 516
rect 11506 572 11570 576
rect 11506 516 11510 572
rect 11510 516 11566 572
rect 11566 516 11570 572
rect 11506 512 11570 516
rect 11586 572 11650 576
rect 11586 516 11590 572
rect 11590 516 11646 572
rect 11646 516 11650 572
rect 11586 512 11650 516
rect 11666 572 11730 576
rect 11666 516 11670 572
rect 11670 516 11726 572
rect 11726 516 11730 572
rect 11666 512 11730 516
rect 11746 572 11810 576
rect 11746 516 11750 572
rect 11750 516 11806 572
rect 11806 516 11810 572
rect 11746 512 11810 516
rect 15208 572 15272 576
rect 15208 516 15212 572
rect 15212 516 15268 572
rect 15268 516 15272 572
rect 15208 512 15272 516
rect 15288 572 15352 576
rect 15288 516 15292 572
rect 15292 516 15348 572
rect 15348 516 15352 572
rect 15288 512 15352 516
rect 15368 572 15432 576
rect 15368 516 15372 572
rect 15372 516 15428 572
rect 15428 516 15432 572
rect 15368 512 15432 516
rect 15448 572 15512 576
rect 15448 516 15452 572
rect 15452 516 15508 572
rect 15508 516 15512 572
rect 15448 512 15512 516
<< metal4 >>
rect 2243 6560 2563 6576
rect 2243 6496 2251 6560
rect 2315 6496 2331 6560
rect 2395 6496 2411 6560
rect 2475 6496 2491 6560
rect 2555 6496 2563 6560
rect 2243 5472 2563 6496
rect 2243 5408 2251 5472
rect 2315 5408 2331 5472
rect 2395 5408 2411 5472
rect 2475 5408 2491 5472
rect 2555 5408 2563 5472
rect 2243 4384 2563 5408
rect 2243 4320 2251 4384
rect 2315 4320 2331 4384
rect 2395 4320 2411 4384
rect 2475 4320 2491 4384
rect 2555 4320 2563 4384
rect 2243 3296 2563 4320
rect 2243 3232 2251 3296
rect 2315 3232 2331 3296
rect 2395 3232 2411 3296
rect 2475 3232 2491 3296
rect 2555 3232 2563 3296
rect 2243 2208 2563 3232
rect 2243 2144 2251 2208
rect 2315 2144 2331 2208
rect 2395 2144 2411 2208
rect 2475 2144 2491 2208
rect 2555 2144 2563 2208
rect 2243 1120 2563 2144
rect 2243 1056 2251 1120
rect 2315 1056 2331 1120
rect 2395 1056 2411 1120
rect 2475 1056 2491 1120
rect 2555 1056 2563 1120
rect 2243 496 2563 1056
rect 4094 6016 4414 6576
rect 4094 5952 4102 6016
rect 4166 5952 4182 6016
rect 4246 5952 4262 6016
rect 4326 5952 4342 6016
rect 4406 5952 4414 6016
rect 4094 4928 4414 5952
rect 4094 4864 4102 4928
rect 4166 4864 4182 4928
rect 4246 4864 4262 4928
rect 4326 4864 4342 4928
rect 4406 4864 4414 4928
rect 4094 3840 4414 4864
rect 4094 3776 4102 3840
rect 4166 3776 4182 3840
rect 4246 3776 4262 3840
rect 4326 3776 4342 3840
rect 4406 3776 4414 3840
rect 4094 2752 4414 3776
rect 4094 2688 4102 2752
rect 4166 2688 4182 2752
rect 4246 2688 4262 2752
rect 4326 2688 4342 2752
rect 4406 2688 4414 2752
rect 4094 1664 4414 2688
rect 4094 1600 4102 1664
rect 4166 1600 4182 1664
rect 4246 1600 4262 1664
rect 4326 1600 4342 1664
rect 4406 1600 4414 1664
rect 4094 576 4414 1600
rect 4094 512 4102 576
rect 4166 512 4182 576
rect 4246 512 4262 576
rect 4326 512 4342 576
rect 4406 512 4414 576
rect 4094 496 4414 512
rect 5945 6560 6265 6576
rect 5945 6496 5953 6560
rect 6017 6496 6033 6560
rect 6097 6496 6113 6560
rect 6177 6496 6193 6560
rect 6257 6496 6265 6560
rect 5945 5472 6265 6496
rect 5945 5408 5953 5472
rect 6017 5408 6033 5472
rect 6097 5408 6113 5472
rect 6177 5408 6193 5472
rect 6257 5408 6265 5472
rect 5945 4384 6265 5408
rect 5945 4320 5953 4384
rect 6017 4320 6033 4384
rect 6097 4320 6113 4384
rect 6177 4320 6193 4384
rect 6257 4320 6265 4384
rect 5945 3296 6265 4320
rect 5945 3232 5953 3296
rect 6017 3232 6033 3296
rect 6097 3232 6113 3296
rect 6177 3232 6193 3296
rect 6257 3232 6265 3296
rect 5945 2208 6265 3232
rect 5945 2144 5953 2208
rect 6017 2144 6033 2208
rect 6097 2144 6113 2208
rect 6177 2144 6193 2208
rect 6257 2144 6265 2208
rect 5945 1120 6265 2144
rect 5945 1056 5953 1120
rect 6017 1056 6033 1120
rect 6097 1056 6113 1120
rect 6177 1056 6193 1120
rect 6257 1056 6265 1120
rect 5945 496 6265 1056
rect 7796 6016 8116 6576
rect 7796 5952 7804 6016
rect 7868 5952 7884 6016
rect 7948 5952 7964 6016
rect 8028 5952 8044 6016
rect 8108 5952 8116 6016
rect 7796 4928 8116 5952
rect 7796 4864 7804 4928
rect 7868 4864 7884 4928
rect 7948 4864 7964 4928
rect 8028 4864 8044 4928
rect 8108 4864 8116 4928
rect 7796 3840 8116 4864
rect 7796 3776 7804 3840
rect 7868 3776 7884 3840
rect 7948 3776 7964 3840
rect 8028 3776 8044 3840
rect 8108 3776 8116 3840
rect 7796 2752 8116 3776
rect 7796 2688 7804 2752
rect 7868 2688 7884 2752
rect 7948 2688 7964 2752
rect 8028 2688 8044 2752
rect 8108 2688 8116 2752
rect 7796 1664 8116 2688
rect 7796 1600 7804 1664
rect 7868 1600 7884 1664
rect 7948 1600 7964 1664
rect 8028 1600 8044 1664
rect 8108 1600 8116 1664
rect 7796 576 8116 1600
rect 7796 512 7804 576
rect 7868 512 7884 576
rect 7948 512 7964 576
rect 8028 512 8044 576
rect 8108 512 8116 576
rect 7796 496 8116 512
rect 9647 6560 9967 6576
rect 9647 6496 9655 6560
rect 9719 6496 9735 6560
rect 9799 6496 9815 6560
rect 9879 6496 9895 6560
rect 9959 6496 9967 6560
rect 9647 5472 9967 6496
rect 9647 5408 9655 5472
rect 9719 5408 9735 5472
rect 9799 5408 9815 5472
rect 9879 5408 9895 5472
rect 9959 5408 9967 5472
rect 9647 4384 9967 5408
rect 9647 4320 9655 4384
rect 9719 4320 9735 4384
rect 9799 4320 9815 4384
rect 9879 4320 9895 4384
rect 9959 4320 9967 4384
rect 9647 3296 9967 4320
rect 9647 3232 9655 3296
rect 9719 3232 9735 3296
rect 9799 3232 9815 3296
rect 9879 3232 9895 3296
rect 9959 3232 9967 3296
rect 9647 2208 9967 3232
rect 9647 2144 9655 2208
rect 9719 2144 9735 2208
rect 9799 2144 9815 2208
rect 9879 2144 9895 2208
rect 9959 2144 9967 2208
rect 9647 1120 9967 2144
rect 9647 1056 9655 1120
rect 9719 1056 9735 1120
rect 9799 1056 9815 1120
rect 9879 1056 9895 1120
rect 9959 1056 9967 1120
rect 9647 496 9967 1056
rect 11498 6016 11818 6576
rect 11498 5952 11506 6016
rect 11570 5952 11586 6016
rect 11650 5952 11666 6016
rect 11730 5952 11746 6016
rect 11810 5952 11818 6016
rect 11498 4928 11818 5952
rect 11498 4864 11506 4928
rect 11570 4864 11586 4928
rect 11650 4864 11666 4928
rect 11730 4864 11746 4928
rect 11810 4864 11818 4928
rect 11498 3840 11818 4864
rect 13349 6560 13669 6576
rect 13349 6496 13357 6560
rect 13421 6496 13437 6560
rect 13501 6496 13517 6560
rect 13581 6496 13597 6560
rect 13661 6496 13669 6560
rect 13349 5472 13669 6496
rect 13349 5408 13357 5472
rect 13421 5408 13437 5472
rect 13501 5408 13517 5472
rect 13581 5408 13597 5472
rect 13661 5408 13669 5472
rect 13123 4588 13189 4589
rect 13123 4524 13124 4588
rect 13188 4524 13189 4588
rect 13123 4523 13189 4524
rect 11498 3776 11506 3840
rect 11570 3776 11586 3840
rect 11650 3776 11666 3840
rect 11730 3776 11746 3840
rect 11810 3776 11818 3840
rect 11498 2752 11818 3776
rect 11498 2688 11506 2752
rect 11570 2688 11586 2752
rect 11650 2688 11666 2752
rect 11730 2688 11746 2752
rect 11810 2688 11818 2752
rect 11498 1664 11818 2688
rect 11498 1600 11506 1664
rect 11570 1600 11586 1664
rect 11650 1600 11666 1664
rect 11730 1600 11746 1664
rect 11810 1600 11818 1664
rect 11498 576 11818 1600
rect 13126 1325 13186 4523
rect 13349 4384 13669 5408
rect 13349 4320 13357 4384
rect 13421 4320 13437 4384
rect 13501 4320 13517 4384
rect 13581 4320 13597 4384
rect 13661 4320 13669 4384
rect 13349 3296 13669 4320
rect 13349 3232 13357 3296
rect 13421 3232 13437 3296
rect 13501 3232 13517 3296
rect 13581 3232 13597 3296
rect 13661 3232 13669 3296
rect 13349 2208 13669 3232
rect 13349 2144 13357 2208
rect 13421 2144 13437 2208
rect 13501 2144 13517 2208
rect 13581 2144 13597 2208
rect 13661 2144 13669 2208
rect 13123 1324 13189 1325
rect 13123 1260 13124 1324
rect 13188 1260 13189 1324
rect 13123 1259 13189 1260
rect 11498 512 11506 576
rect 11570 512 11586 576
rect 11650 512 11666 576
rect 11730 512 11746 576
rect 11810 512 11818 576
rect 11498 496 11818 512
rect 13349 1120 13669 2144
rect 13349 1056 13357 1120
rect 13421 1056 13437 1120
rect 13501 1056 13517 1120
rect 13581 1056 13597 1120
rect 13661 1056 13669 1120
rect 13349 496 13669 1056
rect 15200 6016 15520 6576
rect 15200 5952 15208 6016
rect 15272 5952 15288 6016
rect 15352 5952 15368 6016
rect 15432 5952 15448 6016
rect 15512 5952 15520 6016
rect 15200 4928 15520 5952
rect 15200 4864 15208 4928
rect 15272 4864 15288 4928
rect 15352 4864 15368 4928
rect 15432 4864 15448 4928
rect 15512 4864 15520 4928
rect 15200 3840 15520 4864
rect 15200 3776 15208 3840
rect 15272 3776 15288 3840
rect 15352 3776 15368 3840
rect 15432 3776 15448 3840
rect 15512 3776 15520 3840
rect 15200 2752 15520 3776
rect 15200 2688 15208 2752
rect 15272 2688 15288 2752
rect 15352 2688 15368 2752
rect 15432 2688 15448 2752
rect 15512 2688 15520 2752
rect 15200 1664 15520 2688
rect 15200 1600 15208 1664
rect 15272 1600 15288 1664
rect 15352 1600 15368 1664
rect 15432 1600 15448 1664
rect 15512 1600 15520 1664
rect 15200 576 15520 1600
rect 15200 512 15208 576
rect 15272 512 15288 576
rect 15352 512 15368 576
rect 15432 512 15448 576
rect 15512 512 15520 576
rect 15200 496 15520 512
use sky130_fd_sc_hd__buf_6  _065_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712769939
transform -1 0 15088 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _066_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712769939
transform 1 0 14168 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _067_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712769939
transform -1 0 14352 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _068_
timestamp 1712769939
transform 1 0 14076 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _069_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712769939
transform 1 0 13984 0 1 4896
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _070_
timestamp 1712769939
transform 1 0 11776 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _071_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712769939
transform -1 0 11684 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _072_
timestamp 1712769939
transform 1 0 13524 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _073_
timestamp 1712769939
transform 1 0 13524 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _074_
timestamp 1712769939
transform 1 0 12512 0 -1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _075_
timestamp 1712769939
transform 1 0 12604 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _076_
timestamp 1712769939
transform -1 0 10764 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _077_
timestamp 1712769939
transform 1 0 10764 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _078_
timestamp 1712769939
transform 1 0 10948 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _079_
timestamp 1712769939
transform -1 0 10856 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _080_
timestamp 1712769939
transform -1 0 13524 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _081_
timestamp 1712769939
transform -1 0 7636 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _082_
timestamp 1712769939
transform -1 0 7544 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _083_
timestamp 1712769939
transform 1 0 9384 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _084_
timestamp 1712769939
transform -1 0 8280 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _085_
timestamp 1712769939
transform -1 0 9200 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _086_
timestamp 1712769939
transform -1 0 9476 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _087_
timestamp 1712769939
transform 1 0 8372 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _088_
timestamp 1712769939
transform -1 0 8464 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _089_
timestamp 1712769939
transform -1 0 5704 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _090_
timestamp 1712769939
transform -1 0 6072 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _091_
timestamp 1712769939
transform 1 0 6532 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _092_
timestamp 1712769939
transform -1 0 6716 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _093_
timestamp 1712769939
transform 1 0 8556 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _094_
timestamp 1712769939
transform -1 0 8556 0 -1 5984
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _095_
timestamp 1712769939
transform 1 0 5428 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _096_
timestamp 1712769939
transform 1 0 5796 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _097_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712769939
transform 1 0 13156 0 -1 3808
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _098_
timestamp 1712769939
transform 1 0 11500 0 1 2720
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _099_
timestamp 1712769939
transform 1 0 13524 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _100_
timestamp 1712769939
transform 1 0 8556 0 1 2720
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _101_
timestamp 1712769939
transform 1 0 6256 0 1 3808
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _102_
timestamp 1712769939
transform -1 0 10672 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _103_
timestamp 1712769939
transform 1 0 12788 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__inv_4  _104_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712769939
transform -1 0 6808 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _105_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712769939
transform -1 0 6256 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _106_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712769939
transform 1 0 4692 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _107_
timestamp 1712769939
transform -1 0 13340 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  _108_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712769939
transform 1 0 14352 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _109_
timestamp 1712769939
transform 1 0 13524 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _110_
timestamp 1712769939
transform -1 0 11500 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _111_
timestamp 1712769939
transform 1 0 12512 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _112_
timestamp 1712769939
transform 1 0 11776 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  _113_
timestamp 1712769939
transform -1 0 11776 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _114_
timestamp 1712769939
transform 1 0 11684 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _115_
timestamp 1712769939
transform 1 0 10948 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  _116_
timestamp 1712769939
transform -1 0 9108 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _117_
timestamp 1712769939
transform 1 0 12236 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _118_
timestamp 1712769939
transform -1 0 12512 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _119_
timestamp 1712769939
transform 1 0 10948 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _120_
timestamp 1712769939
transform -1 0 9660 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _121_
timestamp 1712769939
transform 1 0 9752 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _122_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712769939
transform -1 0 7912 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _123_
timestamp 1712769939
transform 1 0 7360 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _124_
timestamp 1712769939
transform -1 0 7452 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _125_
timestamp 1712769939
transform -1 0 6808 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _126_
timestamp 1712769939
transform -1 0 6900 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _127_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712769939
transform 1 0 5060 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _128_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712769939
transform 1 0 4416 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _129_
timestamp 1712769939
transform 1 0 5796 0 1 544
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _130_
timestamp 1712769939
transform 1 0 6164 0 -1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _131_
timestamp 1712769939
transform 1 0 6164 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _132_
timestamp 1712769939
transform -1 0 10764 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _133_
timestamp 1712769939
transform 1 0 8004 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _134_
timestamp 1712769939
transform -1 0 9476 0 1 544
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _135_
timestamp 1712769939
transform 1 0 6992 0 -1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _136_
timestamp 1712769939
transform -1 0 6164 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _137_
timestamp 1712769939
transform 1 0 2576 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _138_
timestamp 1712769939
transform -1 0 3864 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _139_
timestamp 1712769939
transform 1 0 3220 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _140_
timestamp 1712769939
transform -1 0 5060 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _141_
timestamp 1712769939
transform 1 0 4784 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _142_
timestamp 1712769939
transform 1 0 1932 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _143_
timestamp 1712769939
transform 1 0 3220 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _144_
timestamp 1712769939
transform 1 0 3864 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _145_
timestamp 1712769939
transform 1 0 4048 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _146_
timestamp 1712769939
transform -1 0 6348 0 1 1632
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _147_
timestamp 1712769939
transform -1 0 5428 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _148_
timestamp 1712769939
transform 1 0 5336 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _149_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712769939
transform -1 0 10580 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _150_
timestamp 1712769939
transform -1 0 10120 0 -1 4896
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _151_
timestamp 1712769939
transform 1 0 4784 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _152_
timestamp 1712769939
transform -1 0 4784 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _153_
timestamp 1712769939
transform -1 0 4324 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _154_
timestamp 1712769939
transform -1 0 4232 0 -1 2720
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _155_
timestamp 1712769939
transform 1 0 3404 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _156_
timestamp 1712769939
transform 1 0 3680 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _157_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712769939
transform -1 0 3128 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _158_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712769939
transform 1 0 2116 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _159_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712769939
transform 1 0 2116 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _160_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712769939
transform 1 0 2852 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_2  _161_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712769939
transform -1 0 4140 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _162_
timestamp 1712769939
transform -1 0 3588 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _163_
timestamp 1712769939
transform 1 0 2576 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _164_
timestamp 1712769939
transform 1 0 2208 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _165_
timestamp 1712769939
transform 1 0 1748 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _166_
timestamp 1712769939
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _167_
timestamp 1712769939
transform 1 0 1012 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _168_
timestamp 1712769939
transform -1 0 1380 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  clone1
timestamp 1712769939
transform 1 0 11776 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  clone2
timestamp 1712769939
transform -1 0 11592 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_3 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712769939
transform 1 0 828 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_7 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712769939
transform 1 0 1196 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_18
timestamp 1712769939
transform 1 0 2208 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_26 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712769939
transform 1 0 2944 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_32 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712769939
transform 1 0 3496 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_36
timestamp 1712769939
transform 1 0 3864 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_40
timestamp 1712769939
transform 1 0 4232 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_51
timestamp 1712769939
transform 1 0 5244 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55
timestamp 1712769939
transform 1 0 5612 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_67 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712769939
transform 1 0 6716 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_73
timestamp 1712769939
transform 1 0 7268 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_85
timestamp 1712769939
transform 1 0 8372 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_89
timestamp 1712769939
transform 1 0 8740 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_100
timestamp 1712769939
transform 1 0 9752 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_106 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712769939
transform 1 0 10304 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_113
timestamp 1712769939
transform 1 0 10948 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_117
timestamp 1712769939
transform 1 0 11316 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_128
timestamp 1712769939
transform 1 0 12328 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 1712769939
transform 1 0 13340 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_153
timestamp 1712769939
transform 1 0 14628 0 1 544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712769939
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_15
timestamp 1712769939
transform 1 0 1932 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_21
timestamp 1712769939
transform 1 0 2484 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_36
timestamp 1712769939
transform 1 0 3864 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_57
timestamp 1712769939
transform 1 0 5796 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_79
timestamp 1712769939
transform 1 0 7820 0 -1 1632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_88
timestamp 1712769939
transform 1 0 8648 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_100
timestamp 1712769939
transform 1 0 9752 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1712769939
transform 1 0 10764 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_113
timestamp 1712769939
transform 1 0 10948 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_121
timestamp 1712769939
transform 1 0 11684 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_129
timestamp 1712769939
transform 1 0 12420 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_147
timestamp 1712769939
transform 1 0 14076 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_156
timestamp 1712769939
transform 1 0 14904 0 -1 1632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1712769939
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1712769939
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1712769939
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_36
timestamp 1712769939
transform 1 0 3864 0 1 1632
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_63
timestamp 1712769939
transform 1 0 6348 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_75
timestamp 1712769939
transform 1 0 7452 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_79
timestamp 1712769939
transform 1 0 7820 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_94
timestamp 1712769939
transform 1 0 9200 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_105
timestamp 1712769939
transform 1 0 10212 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_135
timestamp 1712769939
transform 1 0 12972 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1712769939
transform 1 0 13340 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_141
timestamp 1712769939
transform 1 0 13524 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_156
timestamp 1712769939
transform 1 0 14904 0 1 1632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1712769939
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_15
timestamp 1712769939
transform 1 0 1932 0 -1 2720
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_40
timestamp 1712769939
transform 1 0 4232 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_52
timestamp 1712769939
transform 1 0 5336 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_57
timestamp 1712769939
transform 1 0 5796 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_67
timestamp 1712769939
transform 1 0 6716 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_79
timestamp 1712769939
transform 1 0 7820 0 -1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_86
timestamp 1712769939
transform 1 0 8464 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_98
timestamp 1712769939
transform 1 0 9568 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_106
timestamp 1712769939
transform 1 0 10304 0 -1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_122
timestamp 1712769939
transform 1 0 11776 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_134
timestamp 1712769939
transform 1 0 12880 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_147
timestamp 1712769939
transform 1 0 14076 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_157
timestamp 1712769939
transform 1 0 14996 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1712769939
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1712769939
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1712769939
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_29
timestamp 1712769939
transform 1 0 3220 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_37
timestamp 1712769939
transform 1 0 3956 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_49
timestamp 1712769939
transform 1 0 5060 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_55
timestamp 1712769939
transform 1 0 5612 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_74
timestamp 1712769939
transform 1 0 7360 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_82
timestamp 1712769939
transform 1 0 8096 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_85
timestamp 1712769939
transform 1 0 8372 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_108
timestamp 1712769939
transform 1 0 10488 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_156
timestamp 1712769939
transform 1 0 14904 0 1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1712769939
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1712769939
transform 1 0 1932 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_27
timestamp 1712769939
transform 1 0 3036 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_40
timestamp 1712769939
transform 1 0 4232 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_44
timestamp 1712769939
transform 1 0 4600 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_53
timestamp 1712769939
transform 1 0 5428 0 -1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_60
timestamp 1712769939
transform 1 0 6072 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_72
timestamp 1712769939
transform 1 0 7176 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_84
timestamp 1712769939
transform 1 0 8280 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_94
timestamp 1712769939
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_107
timestamp 1712769939
transform 1 0 10396 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1712769939
transform 1 0 10764 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_113
timestamp 1712769939
transform 1 0 10948 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_119
timestamp 1712769939
transform 1 0 11500 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_131
timestamp 1712769939
transform 1 0 12604 0 -1 3808
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1712769939
transform 1 0 828 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_22
timestamp 1712769939
transform 1 0 2576 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_41
timestamp 1712769939
transform 1 0 4324 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1712769939
transform 1 0 8188 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_97
timestamp 1712769939
transform 1 0 9476 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_119
timestamp 1712769939
transform 1 0 11500 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1712769939
transform 1 0 13340 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_150
timestamp 1712769939
transform 1 0 14352 0 1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1712769939
transform 1 0 828 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_15
timestamp 1712769939
transform 1 0 1932 0 -1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_23
timestamp 1712769939
transform 1 0 2668 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_35
timestamp 1712769939
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1712769939
transform 1 0 5244 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1712769939
transform 1 0 5612 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_62
timestamp 1712769939
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_109
timestamp 1712769939
transform 1 0 10580 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_131
timestamp 1712769939
transform 1 0 12604 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_142
timestamp 1712769939
transform 1 0 13616 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_147
timestamp 1712769939
transform 1 0 14076 0 -1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1712769939
transform 1 0 828 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_15
timestamp 1712769939
transform 1 0 1932 0 1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1712769939
transform 1 0 3220 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_41
timestamp 1712769939
transform 1 0 4324 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_45
timestamp 1712769939
transform 1 0 4692 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_55
timestamp 1712769939
transform 1 0 5612 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_60
timestamp 1712769939
transform 1 0 6072 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_68
timestamp 1712769939
transform 1 0 6808 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_76
timestamp 1712769939
transform 1 0 7544 0 1 4896
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1712769939
transform 1 0 8372 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_97
timestamp 1712769939
transform 1 0 9476 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_101
timestamp 1712769939
transform 1 0 9844 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_114
timestamp 1712769939
transform 1 0 11040 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_126
timestamp 1712769939
transform 1 0 12144 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1712769939
transform 1 0 13340 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_145
timestamp 1712769939
transform 1 0 13892 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_156
timestamp 1712769939
transform 1 0 14904 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_3
timestamp 1712769939
transform 1 0 828 0 -1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_13
timestamp 1712769939
transform 1 0 1748 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_39
timestamp 1712769939
transform 1 0 4140 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_57
timestamp 1712769939
transform 1 0 5796 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_96
timestamp 1712769939
transform 1 0 9384 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_131
timestamp 1712769939
transform 1 0 12604 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_156
timestamp 1712769939
transform 1 0 14904 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_3
timestamp 1712769939
transform 1 0 828 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_11
timestamp 1712769939
transform 1 0 1564 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_17
timestamp 1712769939
transform 1 0 2116 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_26
timestamp 1712769939
transform 1 0 2944 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_33
timestamp 1712769939
transform 1 0 3588 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_69
timestamp 1712769939
transform 1 0 6900 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_75
timestamp 1712769939
transform 1 0 7452 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_80
timestamp 1712769939
transform 1 0 7912 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_85
timestamp 1712769939
transform 1 0 8372 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_102
timestamp 1712769939
transform 1 0 9936 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_106
timestamp 1712769939
transform 1 0 10304 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_110
timestamp 1712769939
transform 1 0 10672 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_122
timestamp 1712769939
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1712769939
transform 1 0 13340 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_141
timestamp 1712769939
transform 1 0 13524 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_156
timestamp 1712769939
transform 1 0 14904 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1712769939
transform -1 0 15088 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1712769939
transform 1 0 4968 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712769939
transform -1 0 4232 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1712769939
transform 1 0 3220 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1712769939
transform 1 0 1932 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1712769939
transform 1 0 920 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1712769939
transform 1 0 14352 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1712769939
transform 1 0 13064 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1712769939
transform -1 0 12328 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1712769939
transform 1 0 11040 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1712769939
transform -1 0 10304 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1712769939
transform 1 0 9476 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1712769939
transform -1 0 8280 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1712769939
transform 1 0 6992 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1712769939
transform -1 0 6716 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input16
timestamp 1712769939
transform -1 0 15088 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1712769939
transform -1 0 14628 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input18
timestamp 1712769939
transform -1 0 14076 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input19
timestamp 1712769939
transform -1 0 14076 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1712769939
transform 1 0 14628 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1712769939
transform 1 0 14352 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1712769939
transform -1 0 14904 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1712769939
transform 1 0 14352 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1712769939
transform 1 0 14628 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input25
timestamp 1712769939
transform -1 0 13340 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1712769939
transform 1 0 11868 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1712769939
transform 1 0 11592 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1712769939
transform 1 0 10580 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input29
timestamp 1712769939
transform -1 0 10672 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1712769939
transform 1 0 10028 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input31
timestamp 1712769939
transform -1 0 9936 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__maj3_2  mg10 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712769939
transform 1 0 13524 0 1 544
box -38 -48 866 592
use sky130_fd_sc_hd__maj3_1  mg11 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712769939
transform -1 0 14076 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__maj3_2  mg12
timestamp 1712769939
transform 1 0 10948 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__maj3_1  mg13
timestamp 1712769939
transform 1 0 7084 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__maj3_2  mg14
timestamp 1712769939
transform 1 0 8372 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__maj3_1  mg15
timestamp 1712769939
transform 1 0 4692 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__maj3_2  mg16
timestamp 1712769939
transform 1 0 5704 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__maj3_4  mg20 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712769939
transform -1 0 14076 0 -1 2720
box -38 -48 1050 592
use sky130_fd_sc_hd__maj3_2  mg21
timestamp 1712769939
transform 1 0 10672 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__maj3_4  mg22
timestamp 1712769939
transform 1 0 9384 0 -1 3808
box -38 -48 1050 592
use sky130_fd_sc_hd__maj3_4  mg30
timestamp 1712769939
transform 1 0 11592 0 -1 3808
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_11
timestamp 1712769939
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1712769939
transform -1 0 15364 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_12
timestamp 1712769939
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1712769939
transform -1 0 15364 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_13
timestamp 1712769939
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1712769939
transform -1 0 15364 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_14
timestamp 1712769939
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1712769939
transform -1 0 15364 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_15
timestamp 1712769939
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1712769939
transform -1 0 15364 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_16
timestamp 1712769939
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1712769939
transform -1 0 15364 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_17
timestamp 1712769939
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1712769939
transform -1 0 15364 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_18
timestamp 1712769939
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1712769939
transform -1 0 15364 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_19
timestamp 1712769939
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1712769939
transform -1 0 15364 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_20
timestamp 1712769939
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1712769939
transform -1 0 15364 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_21
timestamp 1712769939
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1712769939
transform -1 0 15364 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_22 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712769939
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_23
timestamp 1712769939
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_24
timestamp 1712769939
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_25
timestamp 1712769939
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_26
timestamp 1712769939
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_27
timestamp 1712769939
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_28
timestamp 1712769939
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_29
timestamp 1712769939
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_30
timestamp 1712769939
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_31
timestamp 1712769939
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_32
timestamp 1712769939
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_33
timestamp 1712769939
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_34
timestamp 1712769939
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_35
timestamp 1712769939
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_36
timestamp 1712769939
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_37
timestamp 1712769939
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_38
timestamp 1712769939
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_39
timestamp 1712769939
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_40
timestamp 1712769939
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_41
timestamp 1712769939
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_42
timestamp 1712769939
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_43
timestamp 1712769939
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_44
timestamp 1712769939
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_45
timestamp 1712769939
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_46
timestamp 1712769939
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_47
timestamp 1712769939
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_48
timestamp 1712769939
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_49
timestamp 1712769939
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_50
timestamp 1712769939
transform 1 0 5704 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_51
timestamp 1712769939
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_52
timestamp 1712769939
transform 1 0 10856 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_53
timestamp 1712769939
transform 1 0 13432 0 1 5984
box -38 -48 130 592
<< labels >>
flabel metal4 s 4094 496 4414 6576 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 7796 496 8116 6576 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 11498 496 11818 6576 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 15200 496 15520 6576 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2243 496 2563 6576 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 5945 496 6265 6576 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 9647 496 9967 6576 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 13349 496 13669 6576 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 15014 0 15070 400 0 FreeSans 224 90 0 0 from_adc[0]
port 2 nsew signal input
flabel metal2 s 4894 0 4950 400 0 FreeSans 224 90 0 0 from_adc[10]
port 3 nsew signal input
flabel metal2 s 3882 0 3938 400 0 FreeSans 224 90 0 0 from_adc[11]
port 4 nsew signal input
flabel metal2 s 2870 0 2926 400 0 FreeSans 224 90 0 0 from_adc[12]
port 5 nsew signal input
flabel metal2 s 1858 0 1914 400 0 FreeSans 224 90 0 0 from_adc[13]
port 6 nsew signal input
flabel metal2 s 846 0 902 400 0 FreeSans 224 90 0 0 from_adc[14]
port 7 nsew signal input
flabel metal2 s 14002 0 14058 400 0 FreeSans 224 90 0 0 from_adc[1]
port 8 nsew signal input
flabel metal2 s 12990 0 13046 400 0 FreeSans 224 90 0 0 from_adc[2]
port 9 nsew signal input
flabel metal2 s 11978 0 12034 400 0 FreeSans 224 90 0 0 from_adc[3]
port 10 nsew signal input
flabel metal2 s 10966 0 11022 400 0 FreeSans 224 90 0 0 from_adc[4]
port 11 nsew signal input
flabel metal2 s 9954 0 10010 400 0 FreeSans 224 90 0 0 from_adc[5]
port 12 nsew signal input
flabel metal2 s 8942 0 8998 400 0 FreeSans 224 90 0 0 from_adc[6]
port 13 nsew signal input
flabel metal2 s 7930 0 7986 400 0 FreeSans 224 90 0 0 from_adc[7]
port 14 nsew signal input
flabel metal2 s 6918 0 6974 400 0 FreeSans 224 90 0 0 from_adc[8]
port 15 nsew signal input
flabel metal2 s 5906 0 5962 400 0 FreeSans 224 90 0 0 from_adc[9]
port 16 nsew signal input
flabel metal2 s 15106 6800 15162 7200 0 FreeSans 224 90 0 0 ui_in[0]
port 17 nsew signal input
flabel metal2 s 14738 6800 14794 7200 0 FreeSans 224 90 0 0 ui_in[1]
port 18 nsew signal input
flabel metal2 s 14370 6800 14426 7200 0 FreeSans 224 90 0 0 ui_in[2]
port 19 nsew signal input
flabel metal2 s 14002 6800 14058 7200 0 FreeSans 224 90 0 0 ui_in[3]
port 20 nsew signal input
flabel metal2 s 13634 6800 13690 7200 0 FreeSans 224 90 0 0 ui_in[4]
port 21 nsew signal input
flabel metal2 s 13266 6800 13322 7200 0 FreeSans 224 90 0 0 ui_in[5]
port 22 nsew signal input
flabel metal2 s 12898 6800 12954 7200 0 FreeSans 224 90 0 0 ui_in[6]
port 23 nsew signal input
flabel metal2 s 12530 6800 12586 7200 0 FreeSans 224 90 0 0 ui_in[7]
port 24 nsew signal input
flabel metal2 s 12162 6800 12218 7200 0 FreeSans 224 90 0 0 uio_in[0]
port 25 nsew signal input
flabel metal2 s 11794 6800 11850 7200 0 FreeSans 224 90 0 0 uio_in[1]
port 26 nsew signal input
flabel metal2 s 11426 6800 11482 7200 0 FreeSans 224 90 0 0 uio_in[2]
port 27 nsew signal input
flabel metal2 s 11058 6800 11114 7200 0 FreeSans 224 90 0 0 uio_in[3]
port 28 nsew signal input
flabel metal2 s 10690 6800 10746 7200 0 FreeSans 224 90 0 0 uio_in[4]
port 29 nsew signal input
flabel metal2 s 10322 6800 10378 7200 0 FreeSans 224 90 0 0 uio_in[5]
port 30 nsew signal input
flabel metal2 s 9954 6800 10010 7200 0 FreeSans 224 90 0 0 uio_in[6]
port 31 nsew signal input
flabel metal2 s 9586 6800 9642 7200 0 FreeSans 224 90 0 0 uio_in[7]
port 32 nsew signal input
flabel metal2 s 3330 6800 3386 7200 0 FreeSans 224 90 0 0 uio_oe[0]
port 33 nsew signal tristate
flabel metal2 s 2962 6800 3018 7200 0 FreeSans 224 90 0 0 uio_oe[1]
port 34 nsew signal tristate
flabel metal2 s 2594 6800 2650 7200 0 FreeSans 224 90 0 0 uio_oe[2]
port 35 nsew signal tristate
flabel metal2 s 2226 6800 2282 7200 0 FreeSans 224 90 0 0 uio_oe[3]
port 36 nsew signal tristate
flabel metal2 s 1858 6800 1914 7200 0 FreeSans 224 90 0 0 uio_oe[4]
port 37 nsew signal tristate
flabel metal2 s 1490 6800 1546 7200 0 FreeSans 224 90 0 0 uio_oe[5]
port 38 nsew signal tristate
flabel metal2 s 1122 6800 1178 7200 0 FreeSans 224 90 0 0 uio_oe[6]
port 39 nsew signal tristate
flabel metal2 s 754 6800 810 7200 0 FreeSans 224 90 0 0 uio_oe[7]
port 40 nsew signal tristate
flabel metal2 s 6274 6800 6330 7200 0 FreeSans 224 90 0 0 uio_out[0]
port 41 nsew signal tristate
flabel metal2 s 5906 6800 5962 7200 0 FreeSans 224 90 0 0 uio_out[1]
port 42 nsew signal tristate
flabel metal2 s 5538 6800 5594 7200 0 FreeSans 224 90 0 0 uio_out[2]
port 43 nsew signal tristate
flabel metal2 s 5170 6800 5226 7200 0 FreeSans 224 90 0 0 uio_out[3]
port 44 nsew signal tristate
flabel metal2 s 4802 6800 4858 7200 0 FreeSans 224 90 0 0 uio_out[4]
port 45 nsew signal tristate
flabel metal2 s 4434 6800 4490 7200 0 FreeSans 224 90 0 0 uio_out[5]
port 46 nsew signal tristate
flabel metal2 s 4066 6800 4122 7200 0 FreeSans 224 90 0 0 uio_out[6]
port 47 nsew signal tristate
flabel metal2 s 3698 6800 3754 7200 0 FreeSans 224 90 0 0 uio_out[7]
port 48 nsew signal tristate
flabel metal2 s 9218 6800 9274 7200 0 FreeSans 224 90 0 0 uo_out[0]
port 49 nsew signal tristate
flabel metal2 s 8850 6800 8906 7200 0 FreeSans 224 90 0 0 uo_out[1]
port 50 nsew signal tristate
flabel metal2 s 8482 6800 8538 7200 0 FreeSans 224 90 0 0 uo_out[2]
port 51 nsew signal tristate
flabel metal2 s 8114 6800 8170 7200 0 FreeSans 224 90 0 0 uo_out[3]
port 52 nsew signal tristate
flabel metal2 s 7746 6800 7802 7200 0 FreeSans 224 90 0 0 uo_out[4]
port 53 nsew signal tristate
flabel metal2 s 7378 6800 7434 7200 0 FreeSans 224 90 0 0 uo_out[5]
port 54 nsew signal tristate
flabel metal2 s 7010 6800 7066 7200 0 FreeSans 224 90 0 0 uo_out[6]
port 55 nsew signal tristate
flabel metal2 s 6642 6800 6698 7200 0 FreeSans 224 90 0 0 uo_out[7]
port 56 nsew signal tristate
rlabel via1 8036 5984 8036 5984 0 VGND
rlabel metal1 7958 6528 7958 6528 0 VPWR
rlabel metal1 5658 3570 5658 3570 0 _000_
rlabel metal1 14490 3706 14490 3706 0 _001_
rlabel metal1 13294 3094 13294 3094 0 _002_
rlabel metal1 13386 3910 13386 3910 0 _003_
rlabel metal1 10350 3162 10350 3162 0 _004_
rlabel metal1 9913 4046 9913 4046 0 _005_
rlabel metal1 10764 4250 10764 4250 0 _006_
rlabel metal2 12834 5270 12834 5270 0 _007_
rlabel metal1 4232 3502 4232 3502 0 _008_
rlabel metal1 6946 1326 6946 1326 0 _009_
rlabel metal1 14398 5780 14398 5780 0 _010_
rlabel metal1 13248 3162 13248 3162 0 _011_
rlabel metal1 13018 4148 13018 4148 0 _012_
rlabel metal2 12282 4097 12282 4097 0 _013_
rlabel metal1 11868 5882 11868 5882 0 _014_
rlabel metal1 11638 4250 11638 4250 0 _015_
rlabel metal1 10534 4794 10534 4794 0 _016_
rlabel metal1 12328 5338 12328 5338 0 _017_
rlabel metal2 10994 6018 10994 6018 0 _018_
rlabel metal1 9338 5610 9338 5610 0 _019_
rlabel metal2 7406 5508 7406 5508 0 _020_
rlabel metal1 6808 5882 6808 5882 0 _021_
rlabel metal1 5842 782 5842 782 0 _022_
rlabel metal1 5842 850 5842 850 0 _023_
rlabel metal1 6486 986 6486 986 0 _024_
rlabel metal1 6256 1530 6256 1530 0 _025_
rlabel metal1 9246 816 9246 816 0 _026_
rlabel metal1 8832 850 8832 850 0 _027_
rlabel metal1 8188 646 8188 646 0 _028_
rlabel metal1 6992 1530 6992 1530 0 _029_
rlabel metal1 3174 1360 3174 1360 0 _030_
rlabel metal1 3312 1326 3312 1326 0 _031_
rlabel metal1 4186 2822 4186 2822 0 _032_
rlabel metal2 5014 4658 5014 4658 0 _033_
rlabel metal1 3358 4148 3358 4148 0 _034_
rlabel metal1 4048 4250 4048 4250 0 _035_
rlabel metal2 3910 5508 3910 5508 0 _036_
rlabel metal1 4692 2074 4692 2074 0 _037_
rlabel metal2 5382 5066 5382 5066 0 _038_
rlabel metal1 10028 4658 10028 4658 0 _039_
rlabel metal1 6762 4726 6762 4726 0 _040_
rlabel metal1 4784 5338 4784 5338 0 _041_
rlabel metal1 3979 2482 3979 2482 0 _042_
rlabel metal1 2714 2618 2714 2618 0 _043_
rlabel metal1 3542 3706 3542 3706 0 _044_
rlabel metal1 2898 5134 2898 5134 0 _045_
rlabel metal1 2254 4658 2254 4658 0 _046_
rlabel metal2 3542 5134 3542 5134 0 _047_
rlabel metal1 3542 5610 3542 5610 0 _048_
rlabel metal1 11362 1938 11362 1938 0 _049_
rlabel metal1 14260 1870 14260 1870 0 _050_
rlabel metal1 14076 5202 14076 5202 0 _051_
rlabel metal1 11730 1462 11730 1462 0 _052_
rlabel metal1 13708 5134 13708 5134 0 _053_
rlabel metal1 12650 1530 12650 1530 0 _054_
rlabel metal1 10764 5134 10764 5134 0 _055_
rlabel metal1 10856 2074 10856 2074 0 _056_
rlabel metal1 7268 5678 7268 5678 0 _057_
rlabel metal1 7498 5134 7498 5134 0 _058_
rlabel metal1 8786 1802 8786 1802 0 _059_
rlabel metal1 9292 4046 9292 4046 0 _060_
rlabel metal2 8326 2655 8326 2655 0 _061_
rlabel metal1 6026 5168 6026 5168 0 _062_
rlabel metal2 6578 2686 6578 2686 0 _063_
rlabel metal1 8556 5678 8556 5678 0 _064_
rlabel metal2 15042 568 15042 568 0 from_adc[0]
rlabel metal2 4922 415 4922 415 0 from_adc[10]
rlabel metal2 3910 415 3910 415 0 from_adc[11]
rlabel metal2 2898 568 2898 568 0 from_adc[12]
rlabel metal2 1886 568 1886 568 0 from_adc[13]
rlabel metal2 874 568 874 568 0 from_adc[14]
rlabel metal2 14030 568 14030 568 0 from_adc[1]
rlabel metal2 13018 415 13018 415 0 from_adc[2]
rlabel metal2 12006 415 12006 415 0 from_adc[3]
rlabel metal2 10994 415 10994 415 0 from_adc[4]
rlabel metal2 9982 415 9982 415 0 from_adc[5]
rlabel metal2 8970 534 8970 534 0 from_adc[6]
rlabel metal2 7958 398 7958 398 0 from_adc[7]
rlabel metal2 6946 415 6946 415 0 from_adc[8]
rlabel metal2 5934 415 5934 415 0 from_adc[9]
rlabel metal2 13846 1700 13846 1700 0 maj_level1\[0\]
rlabel metal1 13340 1530 13340 1530 0 maj_level1\[1\]
rlabel metal1 13248 2278 13248 2278 0 maj_level1\[2\]
rlabel metal1 9384 2414 9384 2414 0 maj_level1\[3\]
rlabel via1 9798 2941 9798 2941 0 maj_level1\[4\]
rlabel via1 9798 3451 9798 3451 0 maj_level1\[5\]
rlabel metal2 7452 4046 7452 4046 0 maj_level1\[6\]
rlabel metal2 14122 3247 14122 3247 0 maj_level2\[0\]
rlabel metal1 11684 3162 11684 3162 0 maj_level2\[1\]
rlabel metal1 12144 3366 12144 3366 0 maj_level2\[2\]
rlabel metal2 12558 3876 12558 3876 0 maj_level3
rlabel metal1 13386 3638 13386 3638 0 net1
rlabel metal1 11316 986 11316 986 0 net10
rlabel metal1 10304 986 10304 986 0 net11
rlabel metal1 8326 4556 8326 4556 0 net12
rlabel metal1 7866 986 7866 986 0 net13
rlabel metal1 9798 1938 9798 1938 0 net14
rlabel metal1 7452 1530 7452 1530 0 net15
rlabel metal1 14812 4658 14812 4658 0 net16
rlabel metal1 6026 4624 6026 4624 0 net17
rlabel metal1 14030 4794 14030 4794 0 net18
rlabel metal1 5336 1938 5336 1938 0 net19
rlabel metal1 5152 986 5152 986 0 net2
rlabel metal2 14674 2159 14674 2159 0 net20
rlabel metal1 14398 1768 14398 1768 0 net21
rlabel metal1 10396 5066 10396 5066 0 net22
rlabel metal1 13248 3026 13248 3026 0 net23
rlabel metal1 15134 2074 15134 2074 0 net24
rlabel metal1 8602 2890 8602 2890 0 net25
rlabel metal2 9430 4029 9430 4029 0 net26
rlabel metal2 8878 4488 8878 4488 0 net27
rlabel metal1 5198 5644 5198 5644 0 net28
rlabel metal1 7774 2958 7774 2958 0 net29
rlabel metal1 4370 986 4370 986 0 net3
rlabel metal1 9568 5882 9568 5882 0 net30
rlabel metal2 7222 4318 7222 4318 0 net31
rlabel metal1 9338 5678 9338 5678 0 net32
rlabel metal1 10350 5712 10350 5712 0 net33
rlabel metal1 4232 3978 4232 3978 0 net4
rlabel metal1 3450 918 3450 918 0 net5
rlabel metal1 2484 3570 2484 3570 0 net6
rlabel metal1 14674 6086 14674 6086 0 net7
rlabel via2 4094 4029 4094 4029 0 net8
rlabel metal1 13294 5066 13294 5066 0 net9
rlabel metal1 15088 4046 15088 4046 0 ui_in[0]
rlabel metal1 14674 1394 14674 1394 0 ui_in[1]
rlabel metal1 14214 4658 14214 4658 0 ui_in[2]
rlabel metal2 14030 6538 14030 6538 0 ui_in[3]
rlabel metal1 14858 1360 14858 1360 0 ui_in[4]
rlabel metal1 14582 1904 14582 1904 0 ui_in[5]
rlabel metal1 15226 2958 15226 2958 0 ui_in[6]
rlabel metal1 14582 2924 14582 2924 0 ui_in[7]
rlabel metal1 14950 1870 14950 1870 0 uio_in[0]
rlabel metal2 12282 5185 12282 5185 0 uio_in[1]
rlabel metal1 12098 5168 12098 5168 0 uio_in[2]
rlabel metal1 11730 5134 11730 5134 0 uio_in[3]
rlabel metal1 10764 5746 10764 5746 0 uio_in[4]
rlabel metal1 10488 6222 10488 6222 0 uio_in[5]
rlabel metal1 10166 6222 10166 6222 0 uio_in[6]
rlabel metal1 9660 6222 9660 6222 0 uio_in[7]
rlabel metal2 3358 6640 3358 6640 0 uio_oe[0]
rlabel metal1 2898 6426 2898 6426 0 uio_oe[1]
rlabel metal1 2530 6426 2530 6426 0 uio_oe[2]
rlabel metal1 2070 6426 2070 6426 0 uio_oe[3]
rlabel metal1 1748 5882 1748 5882 0 uio_oe[4]
rlabel metal1 1472 6426 1472 6426 0 uio_oe[5]
rlabel metal2 1150 6368 1150 6368 0 uio_oe[6]
rlabel metal1 966 6222 966 6222 0 uio_oe[7]
rlabel metal1 6348 6426 6348 6426 0 uio_out[0]
rlabel metal1 5888 6426 5888 6426 0 uio_out[1]
rlabel metal1 5336 6426 5336 6426 0 uio_out[2]
rlabel metal1 4278 6324 4278 6324 0 uio_out[3]
rlabel metal1 5198 6358 5198 6358 0 uio_out[4]
rlabel metal1 4508 6426 4508 6426 0 uio_out[5]
rlabel metal1 4002 6426 4002 6426 0 uio_out[6]
rlabel metal1 3864 5882 3864 5882 0 uio_out[7]
rlabel metal1 13754 2006 13754 2006 0 unary_input\[0\]
rlabel metal1 8326 2482 8326 2482 0 unary_input\[10\]
rlabel metal1 3358 4046 3358 4046 0 unary_input\[11\]
rlabel metal2 5382 1666 5382 1666 0 unary_input\[12\]
rlabel metal1 6118 2924 6118 2924 0 unary_input\[13\]
rlabel metal2 5842 3162 5842 3162 0 unary_input\[14\]
rlabel metal1 13938 748 13938 748 0 unary_input\[1\]
rlabel metal1 14030 850 14030 850 0 unary_input\[2\]
rlabel via2 2530 4573 2530 4573 0 unary_input\[3\]
rlabel metal1 13340 1462 13340 1462 0 unary_input\[4\]
rlabel metal1 11362 2516 11362 2516 0 unary_input\[5\]
rlabel metal1 10810 2346 10810 2346 0 unary_input\[6\]
rlabel metal1 7268 5066 7268 5066 0 unary_input\[7\]
rlabel via1 5277 1870 5277 1870 0 unary_input\[8\]
rlabel metal1 8740 1870 8740 1870 0 unary_input\[9\]
rlabel metal2 14582 4845 14582 4845 0 uo_out[0]
rlabel metal1 9982 6290 9982 6290 0 uo_out[1]
rlabel metal1 8648 6290 8648 6290 0 uo_out[2]
rlabel metal1 12052 6426 12052 6426 0 uo_out[3]
rlabel metal1 8510 6426 8510 6426 0 uo_out[4]
rlabel metal1 7544 6426 7544 6426 0 uo_out[5]
rlabel metal1 7130 6426 7130 6426 0 uo_out[6]
rlabel metal2 6670 6640 6670 6640 0 uo_out[7]
<< properties >>
string FIXED_BBOX 0 0 16000 7200
<< end >>
