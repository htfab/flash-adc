VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_htfab_flash_adc
  CLASS BLOCK ;
  FOREIGN tt_um_htfab_flash_adc ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 48.000000 ;
    PORT
      LAYER li1 ;
        RECT 45.860 57.700 46.860 57.870 ;
        RECT 68.520 57.700 69.520 57.870 ;
        RECT 91.180 57.700 92.180 57.870 ;
        RECT 113.840 57.700 114.840 57.870 ;
        RECT 45.860 55.150 46.860 55.320 ;
        RECT 68.520 55.150 69.520 55.320 ;
        RECT 91.180 55.150 92.180 55.320 ;
        RECT 113.840 55.150 114.840 55.320 ;
        RECT 45.860 54.610 46.860 54.780 ;
        RECT 68.520 54.610 69.520 54.780 ;
        RECT 91.180 54.610 92.180 54.780 ;
        RECT 113.840 54.610 114.840 54.780 ;
        RECT 45.860 52.060 46.860 52.230 ;
        RECT 68.520 52.060 69.520 52.230 ;
        RECT 91.180 52.060 92.180 52.230 ;
        RECT 113.840 52.060 114.840 52.230 ;
        RECT 42.100 51.505 43.100 51.675 ;
        RECT 64.760 51.505 65.760 51.675 ;
        RECT 87.420 51.505 88.420 51.675 ;
        RECT 110.080 51.505 111.080 51.675 ;
        RECT 42.100 46.865 43.100 47.035 ;
        RECT 64.760 46.865 65.760 47.035 ;
        RECT 87.420 46.865 88.420 47.035 ;
        RECT 110.080 46.865 111.080 47.035 ;
        RECT 42.100 46.325 43.100 46.495 ;
        RECT 64.760 46.325 65.760 46.495 ;
        RECT 87.420 46.325 88.420 46.495 ;
        RECT 110.080 46.325 111.080 46.495 ;
        RECT 42.100 41.685 43.100 41.855 ;
        RECT 64.760 41.685 65.760 41.855 ;
        RECT 87.420 41.685 88.420 41.855 ;
        RECT 110.080 41.685 111.080 41.855 ;
      LAYER mcon ;
        RECT 45.940 57.700 46.780 57.870 ;
        RECT 68.600 57.700 69.440 57.870 ;
        RECT 91.260 57.700 92.100 57.870 ;
        RECT 113.920 57.700 114.760 57.870 ;
        RECT 45.940 55.150 46.780 55.320 ;
        RECT 68.600 55.150 69.440 55.320 ;
        RECT 91.260 55.150 92.100 55.320 ;
        RECT 113.920 55.150 114.760 55.320 ;
        RECT 45.940 54.610 46.780 54.780 ;
        RECT 68.600 54.610 69.440 54.780 ;
        RECT 91.260 54.610 92.100 54.780 ;
        RECT 113.920 54.610 114.760 54.780 ;
        RECT 45.940 52.060 46.780 52.230 ;
        RECT 68.600 52.060 69.440 52.230 ;
        RECT 91.260 52.060 92.100 52.230 ;
        RECT 113.920 52.060 114.760 52.230 ;
        RECT 42.180 51.505 43.020 51.675 ;
        RECT 64.840 51.505 65.680 51.675 ;
        RECT 87.500 51.505 88.340 51.675 ;
        RECT 110.160 51.505 111.000 51.675 ;
        RECT 42.180 46.865 43.020 47.035 ;
        RECT 64.840 46.865 65.680 47.035 ;
        RECT 87.500 46.865 88.340 47.035 ;
        RECT 110.160 46.865 111.000 47.035 ;
        RECT 42.180 46.325 43.020 46.495 ;
        RECT 64.840 46.325 65.680 46.495 ;
        RECT 87.500 46.325 88.340 46.495 ;
        RECT 110.160 46.325 111.000 46.495 ;
        RECT 42.180 41.685 43.020 41.855 ;
        RECT 64.840 41.685 65.680 41.855 ;
        RECT 87.500 41.685 88.340 41.855 ;
        RECT 110.160 41.685 111.000 41.855 ;
      LAYER met1 ;
        RECT 45.880 57.670 46.840 57.900 ;
        RECT 68.540 57.670 69.500 57.900 ;
        RECT 91.200 57.670 92.160 57.900 ;
        RECT 113.860 57.670 114.820 57.900 ;
        RECT 46.265 55.350 46.455 57.670 ;
        RECT 68.925 55.350 69.115 57.670 ;
        RECT 91.585 55.350 91.775 57.670 ;
        RECT 114.245 55.350 114.435 57.670 ;
        RECT 45.880 54.580 46.840 55.350 ;
        RECT 68.540 54.580 69.500 55.350 ;
        RECT 91.200 54.580 92.160 55.350 ;
        RECT 113.860 54.580 114.820 55.350 ;
        RECT 46.265 52.260 46.455 54.580 ;
        RECT 68.925 52.260 69.115 54.580 ;
        RECT 91.585 52.260 91.775 54.580 ;
        RECT 114.245 52.260 114.435 54.580 ;
        RECT 45.880 52.030 46.840 52.260 ;
        RECT 68.540 52.030 69.500 52.260 ;
        RECT 91.200 52.030 92.160 52.260 ;
        RECT 113.860 52.030 114.820 52.260 ;
        RECT 42.120 51.475 43.080 51.705 ;
        RECT 64.780 51.475 65.740 51.705 ;
        RECT 87.440 51.475 88.400 51.705 ;
        RECT 110.100 51.475 111.060 51.705 ;
        RECT 42.505 47.065 42.695 51.475 ;
        RECT 65.165 47.065 65.355 51.475 ;
        RECT 87.825 47.065 88.015 51.475 ;
        RECT 110.485 47.065 110.675 51.475 ;
        RECT 42.120 46.835 43.080 47.065 ;
        RECT 64.780 46.835 65.740 47.065 ;
        RECT 87.440 46.835 88.400 47.065 ;
        RECT 110.100 46.835 111.060 47.065 ;
        RECT 42.130 46.525 43.070 46.835 ;
        RECT 64.790 46.525 65.730 46.835 ;
        RECT 87.450 46.525 88.390 46.835 ;
        RECT 110.110 46.525 111.050 46.835 ;
        RECT 42.120 46.295 43.080 46.525 ;
        RECT 64.780 46.295 65.740 46.525 ;
        RECT 87.440 46.295 88.400 46.525 ;
        RECT 110.100 46.295 111.060 46.525 ;
        RECT 42.505 41.885 42.695 46.295 ;
        RECT 65.165 41.885 65.355 46.295 ;
        RECT 87.825 41.885 88.015 46.295 ;
        RECT 110.485 41.885 110.675 46.295 ;
        RECT 42.120 41.655 43.080 41.885 ;
        RECT 64.780 41.655 65.740 41.885 ;
        RECT 87.440 41.655 88.400 41.885 ;
        RECT 110.100 41.655 111.060 41.885 ;
      LAYER via ;
        RECT 45.940 54.610 46.780 55.320 ;
        RECT 68.600 54.610 69.440 55.320 ;
        RECT 91.260 54.610 92.100 55.320 ;
        RECT 113.920 54.610 114.760 55.320 ;
        RECT 42.180 46.325 43.020 47.035 ;
        RECT 64.840 46.325 65.680 47.035 ;
        RECT 87.500 46.325 88.340 47.035 ;
        RECT 110.160 46.325 111.000 47.035 ;
      LAYER met2 ;
        RECT 45.880 54.580 46.840 55.350 ;
        RECT 68.540 54.580 69.500 55.350 ;
        RECT 91.200 54.580 92.160 55.350 ;
        RECT 113.860 54.580 114.820 55.350 ;
        RECT 46.250 52.000 46.490 54.580 ;
        RECT 53.230 53.650 55.900 54.140 ;
        RECT 49.430 53.410 55.900 53.650 ;
        RECT 49.430 52.000 49.670 53.410 ;
        RECT 53.230 53.140 55.900 53.410 ;
        RECT 46.250 51.760 49.670 52.000 ;
        RECT 46.250 48.960 46.490 51.760 ;
        RECT 42.480 48.720 46.490 48.960 ;
        RECT 42.480 47.060 42.720 48.720 ;
        RECT 42.130 46.300 43.070 47.060 ;
        RECT 54.900 39.375 55.900 53.140 ;
        RECT 68.910 52.000 69.150 54.580 ;
        RECT 75.890 53.650 78.560 54.140 ;
        RECT 72.090 53.410 78.560 53.650 ;
        RECT 72.090 52.000 72.330 53.410 ;
        RECT 75.890 53.140 78.560 53.410 ;
        RECT 68.910 51.760 72.330 52.000 ;
        RECT 68.910 48.960 69.150 51.760 ;
        RECT 65.140 48.720 69.150 48.960 ;
        RECT 65.140 47.060 65.380 48.720 ;
        RECT 64.790 46.300 65.730 47.060 ;
        RECT 77.560 39.375 78.560 53.140 ;
        RECT 91.570 52.000 91.810 54.580 ;
        RECT 98.550 53.650 101.220 54.140 ;
        RECT 94.750 53.410 101.220 53.650 ;
        RECT 94.750 52.000 94.990 53.410 ;
        RECT 98.550 53.140 101.220 53.410 ;
        RECT 91.570 51.760 94.990 52.000 ;
        RECT 91.570 48.960 91.810 51.760 ;
        RECT 87.800 48.720 91.810 48.960 ;
        RECT 87.800 47.060 88.040 48.720 ;
        RECT 87.450 46.300 88.390 47.060 ;
        RECT 100.220 39.375 101.220 53.140 ;
        RECT 114.230 52.000 114.470 54.580 ;
        RECT 121.210 53.650 123.880 54.140 ;
        RECT 117.410 53.410 123.880 53.650 ;
        RECT 117.410 52.000 117.650 53.410 ;
        RECT 121.210 53.140 123.880 53.410 ;
        RECT 114.230 51.760 117.650 52.000 ;
        RECT 114.230 48.960 114.470 51.760 ;
        RECT 110.460 48.720 114.470 48.960 ;
        RECT 110.460 47.060 110.700 48.720 ;
        RECT 110.110 46.300 111.050 47.060 ;
        RECT 122.880 40.420 123.880 53.140 ;
        RECT 122.835 39.420 123.925 40.420 ;
      LAYER via2 ;
        RECT 54.900 39.420 55.900 40.420 ;
        RECT 77.560 39.420 78.560 40.420 ;
        RECT 100.220 39.420 101.220 40.420 ;
        RECT 122.880 39.420 123.880 40.420 ;
      LAYER met3 ;
        RECT 54.875 40.420 55.925 40.445 ;
        RECT 77.535 40.420 78.585 40.445 ;
        RECT 100.195 40.420 101.245 40.445 ;
        RECT 122.855 40.420 123.905 40.445 ;
        RECT 127.850 40.420 128.840 40.450 ;
        RECT 30.880 39.420 128.875 40.420 ;
        RECT 54.875 39.395 55.925 39.420 ;
        RECT 77.535 39.395 78.585 39.420 ;
        RECT 100.195 39.395 101.245 39.420 ;
        RECT 122.855 39.395 123.905 39.420 ;
        RECT 127.850 39.390 128.840 39.420 ;
      LAYER via3 ;
        RECT 127.840 39.420 128.845 40.420 ;
      LAYER met4 ;
        RECT 127.835 40.420 128.850 40.425 ;
        RECT 127.835 39.420 157.350 40.420 ;
        RECT 127.835 39.415 128.850 39.420 ;
        RECT 156.350 0.000 157.350 39.420 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 113.990 174.065 114.370 174.305 ;
      LAYER mcon ;
        RECT 114.145 174.095 114.315 174.265 ;
      LAYER met1 ;
        RECT 114.085 174.250 114.375 174.295 ;
        RECT 114.530 174.250 114.850 174.310 ;
        RECT 114.085 174.110 114.850 174.250 ;
        RECT 114.085 174.065 114.375 174.110 ;
        RECT 114.530 174.050 114.850 174.110 ;
      LAYER via ;
        RECT 114.560 174.050 114.820 174.310 ;
      LAYER met2 ;
        RECT 114.540 189.615 114.840 190.005 ;
        RECT 114.550 187.950 114.830 189.615 ;
        RECT 114.620 174.340 114.760 187.950 ;
        RECT 114.560 174.020 114.820 174.340 ;
      LAYER via2 ;
        RECT 114.540 189.660 114.840 189.960 ;
      LAYER met3 ;
        RECT 147.410 224.760 147.910 225.760 ;
        RECT 147.510 190.950 147.810 224.760 ;
        RECT 114.540 190.650 147.810 190.950 ;
        RECT 114.540 190.190 114.840 190.650 ;
        RECT 114.340 189.430 115.040 190.190 ;
      LAYER via3 ;
        RECT 147.460 224.810 147.860 225.710 ;
      LAYER met4 ;
        RECT 147.410 224.760 147.910 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER li1 ;
        RECT 111.715 160.755 112.055 161.125 ;
      LAYER mcon ;
        RECT 111.845 160.835 112.015 161.005 ;
      LAYER met1 ;
        RECT 112.690 161.470 113.010 161.730 ;
        RECT 111.785 160.990 112.075 161.035 ;
        RECT 112.780 160.990 112.920 161.470 ;
        RECT 111.785 160.850 112.920 160.990 ;
        RECT 111.785 160.805 112.075 160.850 ;
      LAYER via ;
        RECT 112.720 161.470 112.980 161.730 ;
      LAYER met2 ;
        RECT 112.700 189.615 113.000 190.005 ;
        RECT 112.710 187.950 112.990 189.615 ;
        RECT 112.780 161.760 112.920 187.950 ;
        RECT 112.720 161.440 112.980 161.760 ;
      LAYER via2 ;
        RECT 112.700 189.660 113.000 189.960 ;
      LAYER met3 ;
        RECT 143.730 224.760 144.230 225.760 ;
        RECT 143.830 191.950 144.130 224.760 ;
        RECT 112.700 191.650 144.130 191.950 ;
        RECT 112.700 190.190 113.000 191.650 ;
        RECT 112.500 189.430 113.200 190.190 ;
      LAYER via3 ;
        RECT 143.780 224.810 144.180 225.710 ;
      LAYER met4 ;
        RECT 143.730 224.760 144.230 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 108.960 177.075 109.315 177.445 ;
      LAYER mcon ;
        RECT 109.085 177.155 109.255 177.325 ;
      LAYER met1 ;
        RECT 109.025 177.310 109.315 177.355 ;
        RECT 110.850 177.310 111.170 177.370 ;
        RECT 109.025 177.170 111.170 177.310 ;
        RECT 109.025 177.125 109.315 177.170 ;
        RECT 110.850 177.110 111.170 177.170 ;
      LAYER via ;
        RECT 110.880 177.110 111.140 177.370 ;
      LAYER met2 ;
        RECT 110.860 189.615 111.160 190.005 ;
        RECT 110.870 187.950 111.150 189.615 ;
        RECT 110.940 177.400 111.080 187.950 ;
        RECT 110.880 177.080 111.140 177.400 ;
      LAYER via2 ;
        RECT 110.860 189.660 111.160 189.960 ;
      LAYER met3 ;
        RECT 140.050 224.760 140.550 225.760 ;
        RECT 140.150 192.950 140.450 224.760 ;
        RECT 110.850 192.650 140.450 192.950 ;
        RECT 110.860 190.190 111.160 192.650 ;
        RECT 110.660 189.430 111.360 190.190 ;
      LAYER via3 ;
        RECT 140.100 224.810 140.500 225.710 ;
      LAYER met4 ;
        RECT 140.050 224.760 140.550 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 108.960 184.855 109.315 185.225 ;
      LAYER mcon ;
        RECT 109.085 184.975 109.255 185.145 ;
      LAYER met1 ;
        RECT 109.010 184.930 109.330 185.190 ;
      LAYER via ;
        RECT 109.040 184.930 109.300 185.190 ;
      LAYER met2 ;
        RECT 109.020 189.615 109.320 190.005 ;
        RECT 109.030 187.950 109.310 189.615 ;
        RECT 109.100 185.220 109.240 187.950 ;
        RECT 109.040 184.900 109.300 185.220 ;
      LAYER via2 ;
        RECT 109.020 189.660 109.320 189.960 ;
      LAYER met3 ;
        RECT 136.370 224.760 136.870 225.760 ;
        RECT 136.470 193.950 136.770 224.760 ;
        RECT 109.020 193.650 136.770 193.950 ;
        RECT 109.020 190.190 109.320 193.650 ;
        RECT 108.820 189.430 109.520 190.190 ;
      LAYER via3 ;
        RECT 136.420 224.810 136.820 225.710 ;
      LAYER met4 ;
        RECT 136.370 224.760 136.870 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER li1 ;
        RECT 113.105 160.755 113.435 161.125 ;
      LAYER mcon ;
        RECT 113.225 160.835 113.395 161.005 ;
      LAYER met1 ;
        RECT 107.630 161.470 107.950 161.730 ;
        RECT 107.720 160.990 107.860 161.470 ;
        RECT 107.720 160.850 111.540 160.990 ;
        RECT 111.400 160.650 111.540 160.850 ;
        RECT 113.165 160.805 113.455 161.035 ;
        RECT 113.240 160.650 113.380 160.805 ;
        RECT 111.400 160.510 113.380 160.650 ;
      LAYER via ;
        RECT 107.660 161.470 107.920 161.730 ;
      LAYER met2 ;
        RECT 107.180 189.615 107.480 190.005 ;
        RECT 107.190 187.950 107.470 189.615 ;
        RECT 107.260 187.170 107.400 187.950 ;
        RECT 107.260 187.030 107.860 187.170 ;
        RECT 107.720 182.240 107.860 187.030 ;
        RECT 107.720 182.100 108.320 182.240 ;
        RECT 108.180 179.010 108.320 182.100 ;
        RECT 107.720 178.870 108.320 179.010 ;
        RECT 107.720 161.760 107.860 178.870 ;
        RECT 107.660 161.440 107.920 161.760 ;
      LAYER via2 ;
        RECT 107.180 189.660 107.480 189.960 ;
      LAYER met3 ;
        RECT 132.690 224.760 133.190 225.760 ;
        RECT 132.790 194.950 133.090 224.760 ;
        RECT 107.180 194.650 133.090 194.950 ;
        RECT 107.180 190.190 107.480 194.650 ;
        RECT 106.980 189.430 107.680 190.190 ;
      LAYER via3 ;
        RECT 132.740 224.810 133.140 225.710 ;
      LAYER met4 ;
        RECT 132.690 224.760 133.190 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER li1 ;
        RECT 111.725 163.095 112.055 163.465 ;
      LAYER mcon ;
        RECT 111.845 163.215 112.015 163.385 ;
      LAYER met1 ;
        RECT 104.870 164.190 105.190 164.450 ;
        RECT 104.960 163.710 105.100 164.190 ;
        RECT 104.960 163.570 112.000 163.710 ;
        RECT 111.860 163.415 112.000 163.570 ;
        RECT 111.785 163.185 112.075 163.415 ;
      LAYER via ;
        RECT 104.900 164.190 105.160 164.450 ;
      LAYER met2 ;
        RECT 105.340 189.615 105.640 190.005 ;
        RECT 105.350 187.950 105.630 189.615 ;
        RECT 105.420 167.280 105.560 187.950 ;
        RECT 104.960 167.140 105.560 167.280 ;
        RECT 104.960 164.480 105.100 167.140 ;
        RECT 104.900 164.160 105.160 164.480 ;
      LAYER via2 ;
        RECT 105.340 189.660 105.640 189.960 ;
      LAYER met3 ;
        RECT 129.010 224.760 129.510 225.760 ;
        RECT 129.110 195.950 129.410 224.760 ;
        RECT 105.340 195.650 129.410 195.950 ;
        RECT 105.340 190.190 105.640 195.650 ;
        RECT 105.140 189.430 105.840 190.190 ;
      LAYER via3 ;
        RECT 129.060 224.810 129.460 225.710 ;
      LAYER met4 ;
        RECT 129.010 224.760 129.510 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER li1 ;
        RECT 113.095 168.535 113.435 168.905 ;
      LAYER mcon ;
        RECT 113.225 168.655 113.395 168.825 ;
      LAYER met1 ;
        RECT 103.490 187.170 103.810 187.230 ;
        RECT 116.830 187.170 117.150 187.230 ;
        RECT 103.490 187.030 117.150 187.170 ;
        RECT 103.490 186.970 103.810 187.030 ;
        RECT 116.830 186.970 117.150 187.030 ;
        RECT 116.830 168.950 117.150 169.210 ;
        RECT 113.165 168.810 113.455 168.855 ;
        RECT 116.920 168.810 117.060 168.950 ;
        RECT 113.165 168.670 117.060 168.810 ;
        RECT 113.165 168.625 113.455 168.670 ;
      LAYER via ;
        RECT 103.520 186.970 103.780 187.230 ;
        RECT 116.860 186.970 117.120 187.230 ;
        RECT 116.860 168.950 117.120 169.210 ;
      LAYER met2 ;
        RECT 103.500 189.615 103.800 190.005 ;
        RECT 103.510 187.950 103.790 189.615 ;
        RECT 103.580 187.260 103.720 187.950 ;
        RECT 103.520 186.940 103.780 187.260 ;
        RECT 116.860 186.940 117.120 187.260 ;
        RECT 116.920 169.240 117.060 186.940 ;
        RECT 116.860 168.920 117.120 169.240 ;
      LAYER via2 ;
        RECT 103.500 189.660 103.800 189.960 ;
      LAYER met3 ;
        RECT 125.330 224.760 125.830 225.760 ;
        RECT 125.430 196.950 125.730 224.760 ;
        RECT 103.500 196.650 125.730 196.950 ;
        RECT 103.500 190.190 103.800 196.650 ;
        RECT 103.300 189.430 104.000 190.190 ;
      LAYER via3 ;
        RECT 125.380 224.810 125.780 225.710 ;
      LAYER met4 ;
        RECT 125.330 224.760 125.830 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER li1 ;
        RECT 111.725 168.535 112.055 168.905 ;
      LAYER mcon ;
        RECT 111.845 168.655 112.015 168.825 ;
      LAYER met1 ;
        RECT 111.785 168.625 112.075 168.855 ;
        RECT 111.860 168.470 112.000 168.625 ;
        RECT 112.230 168.470 112.550 168.530 ;
        RECT 111.860 168.330 112.550 168.470 ;
        RECT 112.230 168.270 112.550 168.330 ;
      LAYER via ;
        RECT 112.260 168.270 112.520 168.530 ;
      LAYER met2 ;
        RECT 101.660 189.615 101.960 190.005 ;
        RECT 101.670 187.950 101.950 189.615 ;
        RECT 101.740 182.920 101.880 187.950 ;
        RECT 101.280 182.780 101.880 182.920 ;
        RECT 101.280 175.440 101.420 182.780 ;
        RECT 101.280 175.300 102.340 175.440 ;
        RECT 102.200 168.755 102.340 175.300 ;
        RECT 102.130 168.385 102.410 168.755 ;
        RECT 112.250 168.385 112.530 168.755 ;
        RECT 112.260 168.240 112.520 168.385 ;
      LAYER via2 ;
        RECT 101.660 189.660 101.960 189.960 ;
        RECT 102.130 168.430 102.410 168.710 ;
        RECT 112.250 168.430 112.530 168.710 ;
      LAYER met3 ;
        RECT 121.650 224.760 122.150 225.760 ;
        RECT 121.750 197.950 122.050 224.760 ;
        RECT 101.660 197.650 122.050 197.950 ;
        RECT 101.660 190.190 101.960 197.650 ;
        RECT 101.460 189.430 102.160 190.190 ;
        RECT 102.105 168.720 102.435 168.735 ;
        RECT 112.225 168.720 112.555 168.735 ;
        RECT 102.105 168.420 112.555 168.720 ;
        RECT 102.105 168.405 102.435 168.420 ;
        RECT 112.225 168.405 112.555 168.420 ;
      LAYER via3 ;
        RECT 121.700 224.810 122.100 225.710 ;
      LAYER met4 ;
        RECT 121.650 224.760 122.150 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER li1 ;
        RECT 113.105 163.095 113.435 163.465 ;
      LAYER mcon ;
        RECT 113.225 163.215 113.395 163.385 ;
      LAYER met1 ;
        RECT 100.270 187.850 100.590 187.910 ;
        RECT 114.070 187.850 114.390 187.910 ;
        RECT 100.270 187.710 114.390 187.850 ;
        RECT 100.270 187.650 100.590 187.710 ;
        RECT 114.070 187.650 114.390 187.710 ;
        RECT 114.070 163.850 114.390 164.110 ;
        RECT 113.165 163.370 113.455 163.415 ;
        RECT 114.160 163.370 114.300 163.850 ;
        RECT 113.165 163.230 114.300 163.370 ;
        RECT 113.165 163.185 113.455 163.230 ;
      LAYER via ;
        RECT 100.300 187.650 100.560 187.910 ;
        RECT 114.100 187.650 114.360 187.910 ;
        RECT 114.100 163.850 114.360 164.110 ;
      LAYER met2 ;
        RECT 99.820 189.615 100.120 190.005 ;
        RECT 99.830 187.950 100.110 189.615 ;
        RECT 99.900 187.680 100.040 187.950 ;
        RECT 100.300 187.680 100.560 187.940 ;
        RECT 99.900 187.620 100.560 187.680 ;
        RECT 114.100 187.620 114.360 187.940 ;
        RECT 99.900 187.540 100.500 187.620 ;
        RECT 114.160 164.140 114.300 187.620 ;
        RECT 114.100 163.820 114.360 164.140 ;
      LAYER via2 ;
        RECT 99.820 189.660 100.120 189.960 ;
      LAYER met3 ;
        RECT 117.970 224.760 118.470 225.760 ;
        RECT 118.070 198.950 118.370 224.760 ;
        RECT 99.820 198.650 118.370 198.950 ;
        RECT 99.820 190.190 100.120 198.650 ;
        RECT 99.620 189.430 100.320 190.190 ;
      LAYER via3 ;
        RECT 118.020 224.810 118.420 225.710 ;
      LAYER met4 ;
        RECT 117.970 224.760 118.470 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER li1 ;
        RECT 105.275 179.415 105.615 179.785 ;
      LAYER mcon ;
        RECT 105.405 179.535 105.575 179.705 ;
      LAYER met1 ;
        RECT 100.270 179.690 100.590 179.750 ;
        RECT 105.345 179.690 105.635 179.735 ;
        RECT 100.270 179.550 105.635 179.690 ;
        RECT 100.270 179.490 100.590 179.550 ;
        RECT 105.345 179.505 105.635 179.550 ;
      LAYER via ;
        RECT 100.300 179.490 100.560 179.750 ;
      LAYER met2 ;
        RECT 97.980 189.615 98.280 190.005 ;
        RECT 97.990 187.950 98.270 189.615 ;
        RECT 98.520 188.220 99.580 188.360 ;
        RECT 98.060 187.680 98.200 187.950 ;
        RECT 98.520 187.680 98.660 188.220 ;
        RECT 98.060 187.540 98.660 187.680 ;
        RECT 99.440 180.200 99.580 188.220 ;
        RECT 99.440 180.060 100.500 180.200 ;
        RECT 100.360 179.780 100.500 180.060 ;
        RECT 100.300 179.460 100.560 179.780 ;
      LAYER via2 ;
        RECT 97.980 189.660 98.280 189.960 ;
      LAYER met3 ;
        RECT 114.290 224.760 114.790 225.760 ;
        RECT 114.390 199.950 114.690 224.760 ;
        RECT 97.980 199.650 114.690 199.950 ;
        RECT 97.980 190.190 98.280 199.650 ;
        RECT 97.780 189.430 98.480 190.190 ;
      LAYER via3 ;
        RECT 114.340 224.810 114.740 225.710 ;
      LAYER met4 ;
        RECT 114.290 224.760 114.790 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER li1 ;
        RECT 99.305 179.415 99.635 179.785 ;
      LAYER mcon ;
        RECT 99.425 179.535 99.595 179.705 ;
      LAYER met1 ;
        RECT 96.590 180.710 96.910 180.770 ;
        RECT 96.590 180.570 98.200 180.710 ;
        RECT 96.590 180.510 96.910 180.570 ;
        RECT 98.060 180.030 98.200 180.570 ;
        RECT 98.060 179.890 99.580 180.030 ;
        RECT 99.440 179.735 99.580 179.890 ;
        RECT 99.365 179.505 99.655 179.735 ;
      LAYER via ;
        RECT 96.620 180.510 96.880 180.770 ;
      LAYER met2 ;
        RECT 96.140 189.615 96.440 190.005 ;
        RECT 96.150 187.950 96.430 189.615 ;
        RECT 96.220 182.920 96.360 187.950 ;
        RECT 96.220 182.780 96.820 182.920 ;
        RECT 96.680 180.800 96.820 182.780 ;
        RECT 96.620 180.480 96.880 180.800 ;
      LAYER via2 ;
        RECT 96.140 189.660 96.440 189.960 ;
      LAYER met3 ;
        RECT 110.610 224.760 111.110 225.760 ;
        RECT 110.710 200.950 111.010 224.760 ;
        RECT 96.140 200.650 111.010 200.950 ;
        RECT 96.140 190.190 96.440 200.650 ;
        RECT 95.940 189.430 96.640 190.190 ;
      LAYER via3 ;
        RECT 110.660 224.810 111.060 225.710 ;
      LAYER met4 ;
        RECT 110.610 224.760 111.110 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER li1 ;
        RECT 97.925 179.415 98.255 179.785 ;
      LAYER mcon ;
        RECT 98.045 179.535 98.215 179.705 ;
      LAYER met1 ;
        RECT 94.290 180.030 94.610 180.090 ;
        RECT 94.290 179.890 97.280 180.030 ;
        RECT 94.290 179.830 94.610 179.890 ;
        RECT 97.140 179.690 97.280 179.890 ;
        RECT 97.985 179.690 98.275 179.735 ;
        RECT 97.140 179.550 98.275 179.690 ;
        RECT 97.985 179.505 98.275 179.550 ;
      LAYER via ;
        RECT 94.320 179.830 94.580 180.090 ;
      LAYER met2 ;
        RECT 94.300 189.615 94.600 190.005 ;
        RECT 94.310 187.950 94.590 189.615 ;
        RECT 94.380 180.120 94.520 187.950 ;
        RECT 94.320 179.800 94.580 180.120 ;
      LAYER via2 ;
        RECT 94.300 189.660 94.600 189.960 ;
      LAYER met3 ;
        RECT 106.930 224.760 107.430 225.760 ;
        RECT 107.030 201.950 107.330 224.760 ;
        RECT 94.300 201.650 107.330 201.950 ;
        RECT 94.300 190.190 94.600 201.650 ;
        RECT 94.100 189.430 94.800 190.190 ;
      LAYER via3 ;
        RECT 106.980 224.810 107.380 225.710 ;
      LAYER met4 ;
        RECT 106.930 224.760 107.430 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER li1 ;
        RECT 92.865 182.515 93.195 182.885 ;
      LAYER mcon ;
        RECT 92.985 182.595 93.155 182.765 ;
      LAYER met1 ;
        RECT 92.450 183.230 92.770 183.490 ;
        RECT 92.540 182.750 92.680 183.230 ;
        RECT 92.925 182.750 93.215 182.795 ;
        RECT 92.540 182.610 93.215 182.750 ;
        RECT 92.925 182.565 93.215 182.610 ;
      LAYER via ;
        RECT 92.480 183.230 92.740 183.490 ;
      LAYER met2 ;
        RECT 92.460 189.615 92.760 190.005 ;
        RECT 92.470 187.950 92.750 189.615 ;
        RECT 92.540 183.520 92.680 187.950 ;
        RECT 92.480 183.200 92.740 183.520 ;
      LAYER via2 ;
        RECT 92.460 189.660 92.760 189.960 ;
      LAYER met3 ;
        RECT 103.250 224.760 103.750 225.760 ;
        RECT 103.350 202.950 103.650 224.760 ;
        RECT 92.460 202.650 103.650 202.950 ;
        RECT 92.460 190.190 92.760 202.650 ;
        RECT 92.260 189.430 92.960 190.190 ;
      LAYER via3 ;
        RECT 103.300 224.810 103.700 225.710 ;
      LAYER met4 ;
        RECT 103.250 224.760 103.750 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER li1 ;
        RECT 91.935 184.855 92.275 185.225 ;
      LAYER mcon ;
        RECT 92.065 184.975 92.235 185.145 ;
      LAYER met1 ;
        RECT 90.610 185.130 90.930 185.190 ;
        RECT 92.005 185.130 92.295 185.175 ;
        RECT 90.610 184.990 92.295 185.130 ;
        RECT 90.610 184.930 90.930 184.990 ;
        RECT 92.005 184.945 92.295 184.990 ;
      LAYER via ;
        RECT 90.640 184.930 90.900 185.190 ;
      LAYER met2 ;
        RECT 90.620 189.615 90.920 190.005 ;
        RECT 90.630 187.950 90.910 189.615 ;
        RECT 90.700 185.220 90.840 187.950 ;
        RECT 90.640 184.900 90.900 185.220 ;
      LAYER via2 ;
        RECT 90.620 189.660 90.920 189.960 ;
      LAYER met3 ;
        RECT 99.570 224.760 100.070 225.760 ;
        RECT 99.670 203.950 99.970 224.760 ;
        RECT 90.620 203.650 99.970 203.950 ;
        RECT 90.620 190.190 90.920 203.650 ;
        RECT 90.420 189.430 91.120 190.190 ;
      LAYER via3 ;
        RECT 99.620 224.810 100.020 225.710 ;
      LAYER met4 ;
        RECT 99.570 224.760 100.070 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER li1 ;
        RECT 90.105 184.855 90.435 185.225 ;
      LAYER mcon ;
        RECT 90.225 184.975 90.395 185.145 ;
      LAYER met1 ;
        RECT 89.230 185.130 89.550 185.190 ;
        RECT 90.165 185.130 90.455 185.175 ;
        RECT 89.230 184.990 90.455 185.130 ;
        RECT 89.230 184.930 89.550 184.990 ;
        RECT 90.165 184.945 90.455 184.990 ;
      LAYER via ;
        RECT 89.260 184.930 89.520 185.190 ;
      LAYER met2 ;
        RECT 88.780 189.615 89.080 190.005 ;
        RECT 88.790 187.950 89.070 189.615 ;
        RECT 88.860 187.680 89.000 187.950 ;
        RECT 88.860 187.540 89.460 187.680 ;
        RECT 89.320 185.220 89.460 187.540 ;
        RECT 89.260 184.900 89.520 185.220 ;
      LAYER via2 ;
        RECT 88.780 189.660 89.080 189.960 ;
      LAYER met3 ;
        RECT 95.890 224.760 96.390 225.760 ;
        RECT 95.990 204.950 96.290 224.760 ;
        RECT 88.780 204.650 96.290 204.950 ;
        RECT 88.780 190.190 89.080 204.650 ;
        RECT 88.580 189.430 89.280 190.190 ;
      LAYER via3 ;
        RECT 95.940 224.810 96.340 225.710 ;
      LAYER met4 ;
        RECT 95.890 224.760 96.390 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER li1 ;
        RECT 88.255 184.855 88.595 185.225 ;
      LAYER mcon ;
        RECT 88.385 184.975 88.555 185.145 ;
      LAYER met1 ;
        RECT 86.010 185.130 86.330 185.190 ;
        RECT 88.325 185.130 88.615 185.175 ;
        RECT 86.010 184.990 88.615 185.130 ;
        RECT 86.010 184.930 86.330 184.990 ;
        RECT 88.325 184.945 88.615 184.990 ;
      LAYER via ;
        RECT 86.040 184.930 86.300 185.190 ;
      LAYER met2 ;
        RECT 86.940 189.615 87.240 190.005 ;
        RECT 86.950 187.950 87.230 189.615 ;
        RECT 87.020 187.000 87.160 187.950 ;
        RECT 86.100 186.860 87.160 187.000 ;
        RECT 86.100 185.220 86.240 186.860 ;
        RECT 86.040 184.900 86.300 185.220 ;
      LAYER via2 ;
        RECT 86.940 189.660 87.240 189.960 ;
      LAYER met3 ;
        RECT 92.210 224.760 92.710 225.760 ;
        RECT 92.310 205.950 92.610 224.760 ;
        RECT 86.940 205.650 92.610 205.950 ;
        RECT 86.940 190.190 87.240 205.650 ;
        RECT 86.740 189.430 87.440 190.190 ;
      LAYER via3 ;
        RECT 92.260 224.810 92.660 225.710 ;
      LAYER met4 ;
        RECT 92.210 224.760 92.710 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 55.645 185.430 55.900 186.335 ;
        RECT 55.645 184.700 55.815 185.430 ;
        RECT 55.645 184.125 55.900 184.700 ;
      LAYER mcon ;
        RECT 55.725 185.995 55.895 186.165 ;
      LAYER met1 ;
        RECT 55.650 185.950 55.970 186.210 ;
      LAYER via ;
        RECT 55.680 185.950 55.940 186.210 ;
      LAYER met2 ;
        RECT 55.660 189.615 55.960 190.005 ;
        RECT 55.670 187.950 55.950 189.615 ;
        RECT 55.740 186.240 55.880 187.950 ;
        RECT 55.680 185.920 55.940 186.240 ;
      LAYER via2 ;
        RECT 55.660 189.660 55.960 189.960 ;
      LAYER met3 ;
        RECT 29.650 224.760 30.150 225.760 ;
        RECT 29.750 197.950 30.050 224.760 ;
        RECT 29.750 197.650 55.960 197.950 ;
        RECT 55.660 190.190 55.960 197.650 ;
        RECT 55.460 189.430 56.160 190.190 ;
      LAYER via3 ;
        RECT 29.700 224.810 30.100 225.710 ;
      LAYER met4 ;
        RECT 29.650 224.760 30.150 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 52.960 185.430 53.215 186.335 ;
        RECT 53.045 184.700 53.215 185.430 ;
        RECT 52.960 184.125 53.215 184.700 ;
      LAYER mcon ;
        RECT 52.965 185.995 53.135 186.165 ;
      LAYER met1 ;
        RECT 52.905 186.150 53.195 186.195 ;
        RECT 53.810 186.150 54.130 186.210 ;
        RECT 52.905 186.010 54.130 186.150 ;
        RECT 52.905 185.965 53.195 186.010 ;
        RECT 53.810 185.950 54.130 186.010 ;
      LAYER via ;
        RECT 53.840 185.950 54.100 186.210 ;
      LAYER met2 ;
        RECT 53.820 189.615 54.120 190.005 ;
        RECT 53.830 187.950 54.110 189.615 ;
        RECT 53.900 186.240 54.040 187.950 ;
        RECT 53.840 185.920 54.100 186.240 ;
      LAYER via2 ;
        RECT 53.820 189.660 54.120 189.960 ;
      LAYER met3 ;
        RECT 25.970 224.760 26.470 225.760 ;
        RECT 26.070 196.950 26.370 224.760 ;
        RECT 26.070 196.650 54.120 196.950 ;
        RECT 53.820 190.190 54.120 196.650 ;
        RECT 53.620 189.430 54.320 190.190 ;
      LAYER via3 ;
        RECT 26.020 224.810 26.420 225.710 ;
      LAYER met4 ;
        RECT 25.970 224.760 26.470 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 51.120 185.430 51.375 186.335 ;
        RECT 51.205 184.700 51.375 185.430 ;
        RECT 51.120 184.125 51.375 184.700 ;
      LAYER mcon ;
        RECT 51.125 185.995 51.295 186.165 ;
      LAYER met1 ;
        RECT 51.065 186.150 51.355 186.195 ;
        RECT 51.970 186.150 52.290 186.210 ;
        RECT 51.065 186.010 52.290 186.150 ;
        RECT 51.065 185.965 51.355 186.010 ;
        RECT 51.970 185.950 52.290 186.010 ;
      LAYER via ;
        RECT 52.000 185.950 52.260 186.210 ;
      LAYER met2 ;
        RECT 51.980 189.615 52.280 190.005 ;
        RECT 51.990 187.950 52.270 189.615 ;
        RECT 52.060 186.240 52.200 187.950 ;
        RECT 52.000 185.920 52.260 186.240 ;
      LAYER via2 ;
        RECT 51.980 189.660 52.280 189.960 ;
      LAYER met3 ;
        RECT 22.290 224.760 22.790 225.760 ;
        RECT 22.390 195.950 22.690 224.760 ;
        RECT 22.390 195.650 52.280 195.950 ;
        RECT 51.980 190.190 52.280 195.650 ;
        RECT 51.780 189.430 52.480 190.190 ;
      LAYER via3 ;
        RECT 22.340 224.810 22.740 225.710 ;
      LAYER met4 ;
        RECT 22.290 224.760 22.790 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 48.820 185.430 49.075 186.335 ;
        RECT 48.905 184.700 49.075 185.430 ;
        RECT 48.820 184.125 49.075 184.700 ;
      LAYER mcon ;
        RECT 48.825 185.995 48.995 186.165 ;
      LAYER met1 ;
        RECT 48.765 186.150 49.055 186.195 ;
        RECT 49.670 186.150 49.990 186.210 ;
        RECT 48.765 186.010 49.990 186.150 ;
        RECT 48.765 185.965 49.055 186.010 ;
        RECT 49.670 185.950 49.990 186.010 ;
      LAYER via ;
        RECT 49.700 185.950 49.960 186.210 ;
      LAYER met2 ;
        RECT 50.140 189.615 50.440 190.005 ;
        RECT 50.150 187.950 50.430 189.615 ;
        RECT 50.220 187.680 50.360 187.950 ;
        RECT 49.760 187.540 50.360 187.680 ;
        RECT 49.760 186.240 49.900 187.540 ;
        RECT 49.700 185.920 49.960 186.240 ;
      LAYER via2 ;
        RECT 50.140 189.660 50.440 189.960 ;
      LAYER met3 ;
        RECT 18.610 224.760 19.110 225.760 ;
        RECT 18.710 194.950 19.010 224.760 ;
        RECT 18.710 194.650 50.440 194.950 ;
        RECT 50.140 190.190 50.440 194.650 ;
        RECT 49.940 189.430 50.640 190.190 ;
      LAYER via3 ;
        RECT 18.660 224.810 19.060 225.710 ;
      LAYER met4 ;
        RECT 18.610 224.760 19.110 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 46.980 183.040 47.235 183.615 ;
        RECT 47.065 182.310 47.235 183.040 ;
        RECT 46.980 181.405 47.235 182.310 ;
      LAYER mcon ;
        RECT 46.985 183.275 47.155 183.445 ;
      LAYER met1 ;
        RECT 46.925 183.430 47.215 183.475 ;
        RECT 48.290 183.430 48.610 183.490 ;
        RECT 46.925 183.290 48.610 183.430 ;
        RECT 46.925 183.245 47.215 183.290 ;
        RECT 48.290 183.230 48.610 183.290 ;
      LAYER via ;
        RECT 48.320 183.230 48.580 183.490 ;
      LAYER met2 ;
        RECT 48.300 189.615 48.600 190.005 ;
        RECT 48.310 187.950 48.590 189.615 ;
        RECT 48.380 183.520 48.520 187.950 ;
        RECT 48.320 183.200 48.580 183.520 ;
      LAYER via2 ;
        RECT 48.300 189.660 48.600 189.960 ;
      LAYER met3 ;
        RECT 14.930 224.760 15.430 225.760 ;
        RECT 15.030 193.950 15.330 224.760 ;
        RECT 15.030 193.650 48.600 193.950 ;
        RECT 48.300 190.190 48.600 193.650 ;
        RECT 48.100 189.430 48.800 190.190 ;
      LAYER via3 ;
        RECT 14.980 224.810 15.380 225.710 ;
      LAYER met4 ;
        RECT 14.930 224.760 15.430 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER li1 ;
        RECT 45.125 185.875 45.385 186.335 ;
        RECT 45.985 185.875 46.245 186.335 ;
        RECT 45.125 185.705 46.245 185.875 ;
        RECT 45.985 185.455 46.245 185.705 ;
        RECT 45.985 185.285 46.740 185.455 ;
        RECT 46.335 184.775 46.740 185.285 ;
        RECT 45.090 184.605 46.740 184.775 ;
        RECT 45.090 184.215 45.385 184.605 ;
        RECT 45.985 184.215 46.245 184.605 ;
      LAYER mcon ;
        RECT 46.065 185.995 46.235 186.165 ;
      LAYER met1 ;
        RECT 46.005 186.150 46.295 186.195 ;
        RECT 46.450 186.150 46.770 186.210 ;
        RECT 46.005 186.010 46.770 186.150 ;
        RECT 46.005 185.965 46.295 186.010 ;
        RECT 46.450 185.950 46.770 186.010 ;
      LAYER via ;
        RECT 46.480 185.950 46.740 186.210 ;
      LAYER met2 ;
        RECT 46.460 189.615 46.760 190.005 ;
        RECT 46.470 187.950 46.750 189.615 ;
        RECT 46.540 186.240 46.680 187.950 ;
        RECT 46.480 185.920 46.740 186.240 ;
      LAYER via2 ;
        RECT 46.460 189.660 46.760 189.960 ;
      LAYER met3 ;
        RECT 11.250 224.760 11.750 225.760 ;
        RECT 11.350 192.950 11.650 224.760 ;
        RECT 11.350 192.650 46.760 192.950 ;
        RECT 46.460 190.190 46.760 192.650 ;
        RECT 46.260 189.430 46.960 190.190 ;
      LAYER via3 ;
        RECT 11.300 224.810 11.700 225.710 ;
      LAYER met4 ;
        RECT 11.250 224.760 11.750 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 44.605 183.040 44.860 183.615 ;
        RECT 44.605 182.310 44.775 183.040 ;
        RECT 44.605 181.405 44.860 182.310 ;
      LAYER mcon ;
        RECT 44.685 183.275 44.855 183.445 ;
      LAYER met1 ;
        RECT 44.610 183.230 44.930 183.490 ;
      LAYER via ;
        RECT 44.640 183.230 44.900 183.490 ;
      LAYER met2 ;
        RECT 44.620 189.615 44.920 190.005 ;
        RECT 44.630 187.950 44.910 189.615 ;
        RECT 44.700 183.520 44.840 187.950 ;
        RECT 44.640 183.200 44.900 183.520 ;
      LAYER via2 ;
        RECT 44.620 189.660 44.920 189.960 ;
      LAYER met3 ;
        RECT 7.570 224.760 8.070 225.760 ;
        RECT 7.670 191.950 7.970 224.760 ;
        RECT 7.670 191.650 44.920 191.950 ;
        RECT 44.620 190.190 44.920 191.650 ;
        RECT 44.420 189.430 45.120 190.190 ;
      LAYER via3 ;
        RECT 7.620 224.810 8.020 225.710 ;
      LAYER met4 ;
        RECT 7.570 224.760 8.070 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.914000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 44.505 184.625 44.855 185.195 ;
        RECT 47.845 184.855 48.200 185.225 ;
        RECT 50.145 184.855 50.500 185.225 ;
        RECT 51.985 184.855 52.340 185.225 ;
        RECT 56.520 184.855 56.875 185.225 ;
        RECT 45.480 182.515 45.835 182.885 ;
        RECT 46.005 182.515 46.360 182.885 ;
        RECT 71.325 180.115 71.655 180.895 ;
        RECT 70.890 180.095 71.655 180.115 ;
        RECT 72.165 180.095 72.495 180.895 ;
        RECT 70.890 179.925 72.495 180.095 ;
        RECT 70.890 179.335 71.155 179.925 ;
        RECT 70.890 179.155 72.495 179.335 ;
        RECT 71.325 178.685 71.655 179.155 ;
        RECT 72.165 178.685 72.495 179.155 ;
        RECT 69.455 177.105 70.215 177.355 ;
        RECT 91.145 177.105 91.820 177.355 ;
        RECT 91.555 176.745 91.820 177.105 ;
        RECT 60.275 174.315 60.540 174.675 ;
        RECT 59.865 174.065 60.540 174.315 ;
      LAYER mcon ;
        RECT 44.685 184.975 44.855 185.145 ;
        RECT 47.905 184.975 48.075 185.145 ;
        RECT 50.205 184.975 50.375 185.145 ;
        RECT 52.045 184.975 52.215 185.145 ;
        RECT 56.645 184.975 56.815 185.145 ;
        RECT 45.605 182.595 45.775 182.765 ;
        RECT 46.065 182.595 46.235 182.765 ;
        RECT 72.285 178.855 72.455 179.025 ;
        RECT 69.985 177.155 70.155 177.325 ;
        RECT 91.605 176.815 91.775 176.985 ;
        RECT 60.325 174.435 60.495 174.605 ;
      LAYER met1 ;
        RECT 42.770 185.130 43.090 185.190 ;
        RECT 44.625 185.130 44.915 185.175 ;
        RECT 45.530 185.130 45.850 185.190 ;
        RECT 47.845 185.130 48.135 185.175 ;
        RECT 50.145 185.130 50.435 185.175 ;
        RECT 51.985 185.130 52.275 185.175 ;
        RECT 56.585 185.130 56.875 185.175 ;
        RECT 42.770 184.990 56.875 185.130 ;
        RECT 42.770 184.930 43.090 184.990 ;
        RECT 44.625 184.945 44.915 184.990 ;
        RECT 45.530 184.930 45.850 184.990 ;
        RECT 47.845 184.945 48.135 184.990 ;
        RECT 50.145 184.945 50.435 184.990 ;
        RECT 51.985 184.945 52.275 184.990 ;
        RECT 56.585 184.945 56.875 184.990 ;
        RECT 56.660 184.790 56.800 184.945 ;
        RECT 61.630 184.930 61.950 185.190 ;
        RECT 61.720 184.790 61.860 184.930 ;
        RECT 56.660 184.650 61.860 184.790 ;
        RECT 45.530 182.750 45.850 182.810 ;
        RECT 46.005 182.750 46.295 182.795 ;
        RECT 45.530 182.610 46.295 182.750 ;
        RECT 45.530 182.550 45.850 182.610 ;
        RECT 46.005 182.565 46.295 182.610 ;
        RECT 69.910 179.010 70.230 179.070 ;
        RECT 72.225 179.010 72.515 179.055 ;
        RECT 86.470 179.010 86.790 179.070 ;
        RECT 69.910 178.870 86.790 179.010 ;
        RECT 69.910 178.810 70.230 178.870 ;
        RECT 72.225 178.825 72.515 178.870 ;
        RECT 86.470 178.810 86.790 178.870 ;
        RECT 69.910 177.110 70.230 177.370 ;
        RECT 91.545 176.785 91.835 177.015 ;
        RECT 60.250 176.630 60.570 176.690 ;
        RECT 61.630 176.630 61.950 176.690 ;
        RECT 69.910 176.630 70.230 176.690 ;
        RECT 60.250 176.490 70.230 176.630 ;
        RECT 60.250 176.430 60.570 176.490 ;
        RECT 61.630 176.430 61.950 176.490 ;
        RECT 69.910 176.430 70.230 176.490 ;
        RECT 86.470 176.630 86.790 176.690 ;
        RECT 91.620 176.630 91.760 176.785 ;
        RECT 86.470 176.490 91.760 176.630 ;
        RECT 86.470 176.430 86.790 176.490 ;
        RECT 60.250 174.390 60.570 174.650 ;
      LAYER via ;
        RECT 42.800 184.930 43.060 185.190 ;
        RECT 45.560 184.930 45.820 185.190 ;
        RECT 61.660 184.930 61.920 185.190 ;
        RECT 45.560 182.550 45.820 182.810 ;
        RECT 69.940 178.810 70.200 179.070 ;
        RECT 86.500 178.810 86.760 179.070 ;
        RECT 69.940 177.110 70.200 177.370 ;
        RECT 60.280 176.430 60.540 176.690 ;
        RECT 61.660 176.430 61.920 176.690 ;
        RECT 69.940 176.430 70.200 176.690 ;
        RECT 86.500 176.430 86.760 176.690 ;
        RECT 60.280 174.390 60.540 174.650 ;
      LAYER met2 ;
        RECT 42.780 189.615 43.080 190.005 ;
        RECT 42.790 187.950 43.070 189.615 ;
        RECT 42.860 185.220 43.000 187.950 ;
        RECT 42.800 184.900 43.060 185.220 ;
        RECT 45.560 184.900 45.820 185.220 ;
        RECT 61.660 184.900 61.920 185.220 ;
        RECT 45.620 182.840 45.760 184.900 ;
        RECT 45.560 182.520 45.820 182.840 ;
        RECT 61.720 176.720 61.860 184.900 ;
        RECT 69.940 178.780 70.200 179.100 ;
        RECT 86.500 178.780 86.760 179.100 ;
        RECT 70.000 177.400 70.140 178.780 ;
        RECT 69.940 177.080 70.200 177.400 ;
        RECT 70.000 176.720 70.140 177.080 ;
        RECT 86.560 176.720 86.700 178.780 ;
        RECT 60.280 176.400 60.540 176.720 ;
        RECT 61.660 176.400 61.920 176.720 ;
        RECT 69.940 176.400 70.200 176.720 ;
        RECT 86.500 176.400 86.760 176.720 ;
        RECT 60.340 174.680 60.480 176.400 ;
        RECT 60.280 174.360 60.540 174.680 ;
      LAYER via2 ;
        RECT 42.780 189.660 43.080 189.960 ;
      LAYER met3 ;
        RECT 3.890 224.760 4.390 225.760 ;
        RECT 3.990 190.950 4.290 224.760 ;
        RECT 3.990 190.650 43.080 190.950 ;
        RECT 42.780 190.190 43.080 190.650 ;
        RECT 42.580 189.430 43.280 190.190 ;
      LAYER via3 ;
        RECT 3.940 224.810 4.340 225.710 ;
      LAYER met4 ;
        RECT 3.890 224.760 4.390 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 70.900 185.430 71.155 186.335 ;
        RECT 70.985 184.700 71.155 185.430 ;
        RECT 70.900 184.125 71.155 184.700 ;
      LAYER mcon ;
        RECT 70.905 185.995 71.075 186.165 ;
      LAYER met1 ;
        RECT 70.370 186.150 70.690 186.210 ;
        RECT 70.845 186.150 71.135 186.195 ;
        RECT 70.370 186.010 71.135 186.150 ;
        RECT 70.370 185.950 70.690 186.010 ;
        RECT 70.845 185.965 71.135 186.010 ;
      LAYER via ;
        RECT 70.400 185.950 70.660 186.210 ;
      LAYER met2 ;
        RECT 70.380 189.615 70.680 190.005 ;
        RECT 70.390 187.950 70.670 189.615 ;
        RECT 70.460 186.240 70.600 187.950 ;
        RECT 70.400 185.920 70.660 186.240 ;
      LAYER via2 ;
        RECT 70.380 189.660 70.680 189.960 ;
      LAYER met3 ;
        RECT 59.090 224.760 59.590 225.760 ;
        RECT 59.190 205.950 59.490 224.760 ;
        RECT 59.190 205.650 70.680 205.950 ;
        RECT 70.380 190.190 70.680 205.650 ;
        RECT 70.180 189.430 70.880 190.190 ;
      LAYER via3 ;
        RECT 59.140 224.810 59.540 225.710 ;
      LAYER met4 ;
        RECT 59.090 224.760 59.590 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 68.525 185.430 68.780 186.335 ;
        RECT 68.525 184.700 68.695 185.430 ;
        RECT 68.525 184.125 68.780 184.700 ;
      LAYER mcon ;
        RECT 68.605 185.995 68.775 186.165 ;
      LAYER met1 ;
        RECT 68.070 186.150 68.390 186.210 ;
        RECT 68.545 186.150 68.835 186.195 ;
        RECT 68.070 186.010 68.835 186.150 ;
        RECT 68.070 185.950 68.390 186.010 ;
        RECT 68.545 185.965 68.835 186.010 ;
      LAYER via ;
        RECT 68.100 185.950 68.360 186.210 ;
      LAYER met2 ;
        RECT 68.540 189.615 68.840 190.005 ;
        RECT 68.550 187.950 68.830 189.615 ;
        RECT 68.620 187.680 68.760 187.950 ;
        RECT 68.160 187.540 68.760 187.680 ;
        RECT 68.160 186.240 68.300 187.540 ;
        RECT 68.100 185.920 68.360 186.240 ;
      LAYER via2 ;
        RECT 68.540 189.660 68.840 189.960 ;
      LAYER met3 ;
        RECT 55.410 224.760 55.910 225.760 ;
        RECT 55.510 204.950 55.810 224.760 ;
        RECT 55.510 204.650 68.840 204.950 ;
        RECT 68.540 190.190 68.840 204.650 ;
        RECT 68.340 189.430 69.040 190.190 ;
      LAYER via3 ;
        RECT 55.460 224.810 55.860 225.710 ;
      LAYER met4 ;
        RECT 55.410 224.760 55.910 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER li1 ;
        RECT 63.985 185.875 64.245 186.335 ;
        RECT 64.845 185.875 65.105 186.335 ;
        RECT 63.985 185.705 65.105 185.875 ;
        RECT 64.845 185.455 65.105 185.705 ;
        RECT 64.845 185.285 65.600 185.455 ;
        RECT 65.195 184.775 65.600 185.285 ;
        RECT 63.950 184.605 65.600 184.775 ;
        RECT 63.950 184.215 64.245 184.605 ;
        RECT 64.845 184.215 65.105 184.605 ;
      LAYER mcon ;
        RECT 64.925 185.995 65.095 186.165 ;
      LAYER met1 ;
        RECT 64.865 186.150 65.155 186.195 ;
        RECT 66.230 186.150 66.550 186.210 ;
        RECT 64.865 186.010 66.550 186.150 ;
        RECT 64.865 185.965 65.155 186.010 ;
        RECT 66.230 185.950 66.550 186.010 ;
      LAYER via ;
        RECT 66.260 185.950 66.520 186.210 ;
      LAYER met2 ;
        RECT 66.700 189.615 67.000 190.005 ;
        RECT 66.710 187.950 66.990 189.615 ;
        RECT 66.780 186.320 66.920 187.950 ;
        RECT 66.320 186.240 66.920 186.320 ;
        RECT 66.260 186.180 66.920 186.240 ;
        RECT 66.260 185.920 66.520 186.180 ;
      LAYER via2 ;
        RECT 66.700 189.660 67.000 189.960 ;
      LAYER met3 ;
        RECT 51.730 224.760 52.230 225.760 ;
        RECT 51.830 203.950 52.130 224.760 ;
        RECT 51.830 203.650 67.000 203.950 ;
        RECT 66.700 190.190 67.000 203.650 ;
        RECT 66.500 189.430 67.200 190.190 ;
      LAYER via3 ;
        RECT 51.780 224.810 52.180 225.710 ;
      LAYER met4 ;
        RECT 51.730 224.760 52.230 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 60.320 185.430 60.575 186.335 ;
        RECT 60.405 184.700 60.575 185.430 ;
        RECT 60.320 184.125 60.575 184.700 ;
      LAYER mcon ;
        RECT 60.325 185.655 60.495 185.825 ;
      LAYER met1 ;
        RECT 60.265 185.625 60.555 185.855 ;
        RECT 60.340 185.470 60.480 185.625 ;
        RECT 64.850 185.470 65.170 185.530 ;
        RECT 60.340 185.330 65.170 185.470 ;
        RECT 64.850 185.270 65.170 185.330 ;
      LAYER via ;
        RECT 64.880 185.270 65.140 185.530 ;
      LAYER met2 ;
        RECT 64.860 189.615 65.160 190.005 ;
        RECT 64.870 187.950 65.150 189.615 ;
        RECT 64.940 185.560 65.080 187.950 ;
        RECT 64.880 185.240 65.140 185.560 ;
      LAYER via2 ;
        RECT 64.860 189.660 65.160 189.960 ;
      LAYER met3 ;
        RECT 48.050 224.760 48.550 225.760 ;
        RECT 48.150 202.950 48.450 224.760 ;
        RECT 48.150 202.650 65.160 202.950 ;
        RECT 64.860 190.190 65.160 202.650 ;
        RECT 64.660 189.430 65.360 190.190 ;
      LAYER via3 ;
        RECT 48.100 224.810 48.500 225.710 ;
      LAYER met4 ;
        RECT 48.050 224.760 48.550 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 66.760 185.430 67.015 186.335 ;
        RECT 66.845 184.700 67.015 185.430 ;
        RECT 66.760 184.125 67.015 184.700 ;
      LAYER mcon ;
        RECT 66.765 185.655 66.935 185.825 ;
      LAYER met1 ;
        RECT 63.010 185.950 63.330 186.210 ;
        RECT 63.100 185.810 63.240 185.950 ;
        RECT 66.705 185.810 66.995 185.855 ;
        RECT 63.100 185.670 66.995 185.810 ;
        RECT 66.705 185.625 66.995 185.670 ;
      LAYER via ;
        RECT 63.040 185.950 63.300 186.210 ;
      LAYER met2 ;
        RECT 63.020 189.615 63.320 190.005 ;
        RECT 63.030 187.950 63.310 189.615 ;
        RECT 63.100 186.240 63.240 187.950 ;
        RECT 63.040 185.920 63.300 186.240 ;
      LAYER via2 ;
        RECT 63.020 189.660 63.320 189.960 ;
      LAYER met3 ;
        RECT 44.370 224.760 44.870 225.760 ;
        RECT 44.470 201.950 44.770 224.760 ;
        RECT 44.470 201.650 63.320 201.950 ;
        RECT 63.020 190.190 63.320 201.650 ;
        RECT 62.820 189.430 63.520 190.190 ;
      LAYER via3 ;
        RECT 44.420 224.810 44.820 225.710 ;
      LAYER met4 ;
        RECT 44.370 224.760 44.870 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 61.625 185.430 61.880 186.335 ;
        RECT 61.625 184.700 61.795 185.430 ;
        RECT 61.625 184.125 61.880 184.700 ;
      LAYER mcon ;
        RECT 61.705 185.995 61.875 186.165 ;
      LAYER met1 ;
        RECT 61.170 186.150 61.490 186.210 ;
        RECT 61.645 186.150 61.935 186.195 ;
        RECT 61.170 186.010 61.935 186.150 ;
        RECT 61.170 185.950 61.490 186.010 ;
        RECT 61.645 185.965 61.935 186.010 ;
      LAYER via ;
        RECT 61.200 185.950 61.460 186.210 ;
      LAYER met2 ;
        RECT 61.180 189.615 61.480 190.005 ;
        RECT 61.190 187.950 61.470 189.615 ;
        RECT 61.260 186.240 61.400 187.950 ;
        RECT 61.200 185.920 61.460 186.240 ;
      LAYER via2 ;
        RECT 61.180 189.660 61.480 189.960 ;
      LAYER met3 ;
        RECT 40.690 224.760 41.190 225.760 ;
        RECT 40.790 200.950 41.090 224.760 ;
        RECT 40.790 200.650 61.480 200.950 ;
        RECT 61.180 190.190 61.480 200.650 ;
        RECT 60.980 189.430 61.680 190.190 ;
      LAYER via3 ;
        RECT 40.740 224.810 41.140 225.710 ;
      LAYER met4 ;
        RECT 40.690 224.760 41.190 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 58.480 185.430 58.735 186.335 ;
        RECT 58.565 184.700 58.735 185.430 ;
        RECT 58.480 184.125 58.735 184.700 ;
      LAYER mcon ;
        RECT 58.485 185.995 58.655 186.165 ;
      LAYER met1 ;
        RECT 58.425 186.150 58.715 186.195 ;
        RECT 59.330 186.150 59.650 186.210 ;
        RECT 58.425 186.010 59.650 186.150 ;
        RECT 58.425 185.965 58.715 186.010 ;
        RECT 59.330 185.950 59.650 186.010 ;
      LAYER via ;
        RECT 59.360 185.950 59.620 186.210 ;
      LAYER met2 ;
        RECT 59.340 189.615 59.640 190.005 ;
        RECT 59.350 187.950 59.630 189.615 ;
        RECT 59.420 186.240 59.560 187.950 ;
        RECT 59.360 185.920 59.620 186.240 ;
      LAYER via2 ;
        RECT 59.340 189.660 59.640 189.960 ;
      LAYER met3 ;
        RECT 37.010 224.760 37.510 225.760 ;
        RECT 37.110 199.950 37.410 224.760 ;
        RECT 37.110 199.650 59.640 199.950 ;
        RECT 59.340 190.190 59.640 199.650 ;
        RECT 59.140 189.430 59.840 190.190 ;
      LAYER via3 ;
        RECT 37.060 224.810 37.460 225.710 ;
      LAYER met4 ;
        RECT 37.010 224.760 37.510 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.453750 ;
    PORT
      LAYER li1 ;
        RECT 58.945 181.405 59.190 183.615 ;
      LAYER mcon ;
        RECT 58.945 183.275 59.115 183.445 ;
      LAYER met1 ;
        RECT 57.490 183.430 57.810 183.490 ;
        RECT 58.885 183.430 59.175 183.475 ;
        RECT 57.490 183.290 59.175 183.430 ;
        RECT 57.490 183.230 57.810 183.290 ;
        RECT 58.885 183.245 59.175 183.290 ;
      LAYER via ;
        RECT 57.520 183.230 57.780 183.490 ;
      LAYER met2 ;
        RECT 57.500 189.615 57.800 190.005 ;
        RECT 57.510 187.950 57.790 189.615 ;
        RECT 57.580 183.520 57.720 187.950 ;
        RECT 57.520 183.200 57.780 183.520 ;
      LAYER via2 ;
        RECT 57.500 189.660 57.800 189.960 ;
      LAYER met3 ;
        RECT 33.330 224.760 33.830 225.760 ;
        RECT 33.430 198.950 33.730 224.760 ;
        RECT 33.430 198.650 57.800 198.950 ;
        RECT 57.500 190.190 57.800 198.650 ;
        RECT 57.300 189.430 58.000 190.190 ;
      LAYER via3 ;
        RECT 33.380 224.810 33.780 225.710 ;
      LAYER met4 ;
        RECT 33.330 224.760 33.830 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 111.795 183.135 111.965 183.615 ;
        RECT 112.635 183.135 112.805 183.615 ;
        RECT 111.795 182.965 112.805 183.135 ;
        RECT 112.310 182.425 112.805 182.965 ;
        RECT 111.795 182.255 112.805 182.425 ;
        RECT 111.795 181.405 111.965 182.255 ;
        RECT 112.635 181.405 112.805 182.255 ;
      LAYER mcon ;
        RECT 111.845 182.255 112.015 182.425 ;
      LAYER met1 ;
        RECT 111.770 182.210 112.090 182.470 ;
      LAYER via ;
        RECT 111.800 182.210 112.060 182.470 ;
      LAYER met2 ;
        RECT 85.100 189.615 85.400 190.005 ;
        RECT 85.110 187.950 85.390 189.615 ;
        RECT 85.180 174.195 85.320 187.950 ;
        RECT 111.800 182.180 112.060 182.500 ;
        RECT 111.860 174.195 112.000 182.180 ;
        RECT 85.110 173.825 85.390 174.195 ;
        RECT 111.790 173.825 112.070 174.195 ;
      LAYER via2 ;
        RECT 85.100 189.660 85.400 189.960 ;
        RECT 85.110 173.870 85.390 174.150 ;
        RECT 111.790 173.870 112.070 174.150 ;
      LAYER met3 ;
        RECT 88.530 224.760 89.030 225.760 ;
        RECT 88.630 206.950 88.930 224.760 ;
        RECT 85.100 206.650 88.930 206.950 ;
        RECT 85.100 190.190 85.400 206.650 ;
        RECT 84.900 189.430 85.600 190.190 ;
        RECT 85.085 174.160 85.415 174.175 ;
        RECT 111.765 174.160 112.095 174.175 ;
        RECT 85.085 173.860 112.095 174.160 ;
        RECT 85.085 173.845 85.415 173.860 ;
        RECT 111.765 173.845 112.095 173.860 ;
      LAYER via3 ;
        RECT 88.580 224.810 88.980 225.710 ;
      LAYER met4 ;
        RECT 88.530 224.760 89.030 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER li1 ;
        RECT 94.355 185.485 94.525 186.335 ;
        RECT 95.195 185.485 95.365 186.335 ;
        RECT 96.035 185.485 96.205 186.335 ;
        RECT 94.355 185.315 96.205 185.485 ;
        RECT 94.355 184.775 95.690 185.315 ;
        RECT 94.355 184.605 96.205 184.775 ;
        RECT 94.355 184.125 94.525 184.605 ;
        RECT 95.195 184.125 95.365 184.605 ;
        RECT 96.035 184.125 96.205 184.605 ;
      LAYER mcon ;
        RECT 94.365 185.315 94.535 185.485 ;
      LAYER met1 ;
        RECT 83.250 185.610 83.570 185.870 ;
        RECT 83.340 185.470 83.480 185.610 ;
        RECT 94.305 185.470 94.595 185.515 ;
        RECT 83.340 185.330 94.595 185.470 ;
        RECT 94.305 185.285 94.595 185.330 ;
      LAYER via ;
        RECT 83.280 185.610 83.540 185.870 ;
      LAYER met2 ;
        RECT 83.260 189.615 83.560 190.005 ;
        RECT 83.270 187.950 83.550 189.615 ;
        RECT 83.340 185.900 83.480 187.950 ;
        RECT 83.280 185.580 83.540 185.900 ;
      LAYER via2 ;
        RECT 83.260 189.660 83.560 189.960 ;
      LAYER met3 ;
        RECT 84.850 224.760 85.350 225.760 ;
        RECT 84.950 207.950 85.250 224.760 ;
        RECT 83.260 207.650 85.250 207.950 ;
        RECT 83.260 190.190 83.560 207.650 ;
        RECT 83.060 189.430 83.760 190.190 ;
      LAYER via3 ;
        RECT 84.900 224.810 85.300 225.710 ;
      LAYER met4 ;
        RECT 84.850 224.760 85.350 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 82.535 185.485 82.705 186.335 ;
        RECT 83.375 185.485 83.545 186.335 ;
        RECT 82.535 185.315 83.545 185.485 ;
        RECT 82.535 184.775 83.030 185.315 ;
        RECT 82.535 184.605 83.545 184.775 ;
        RECT 82.535 184.125 82.705 184.605 ;
        RECT 83.375 184.125 83.545 184.605 ;
      LAYER mcon ;
        RECT 82.865 185.315 83.035 185.485 ;
      LAYER met1 ;
        RECT 81.410 185.470 81.730 185.530 ;
        RECT 82.805 185.470 83.095 185.515 ;
        RECT 81.410 185.330 83.095 185.470 ;
        RECT 81.410 185.270 81.730 185.330 ;
        RECT 82.805 185.285 83.095 185.330 ;
      LAYER via ;
        RECT 81.440 185.270 81.700 185.530 ;
      LAYER met2 ;
        RECT 81.420 189.615 81.720 190.005 ;
        RECT 81.430 187.950 81.710 189.615 ;
        RECT 81.500 185.560 81.640 187.950 ;
        RECT 81.440 185.240 81.700 185.560 ;
      LAYER via2 ;
        RECT 81.420 189.660 81.720 189.960 ;
      LAYER met3 ;
        RECT 81.170 224.760 81.670 225.760 ;
        RECT 81.270 190.950 81.570 224.760 ;
        RECT 81.270 190.650 81.720 190.950 ;
        RECT 81.420 190.190 81.720 190.650 ;
        RECT 81.220 189.430 81.920 190.190 ;
      LAYER via3 ;
        RECT 81.220 224.810 81.620 225.710 ;
      LAYER met4 ;
        RECT 81.170 224.760 81.670 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER li1 ;
        RECT 99.415 185.875 99.675 186.335 ;
        RECT 100.275 185.875 100.535 186.335 ;
        RECT 99.415 185.705 100.535 185.875 ;
        RECT 99.415 185.455 99.675 185.705 ;
        RECT 98.920 185.285 99.675 185.455 ;
        RECT 98.920 184.775 99.325 185.285 ;
        RECT 98.920 184.605 100.570 184.775 ;
        RECT 99.415 184.215 99.675 184.605 ;
        RECT 100.275 184.215 100.570 184.605 ;
      LAYER mcon ;
        RECT 99.425 185.995 99.595 186.165 ;
      LAYER met1 ;
        RECT 79.570 187.170 79.890 187.230 ;
        RECT 98.890 187.170 99.210 187.230 ;
        RECT 79.570 187.030 99.210 187.170 ;
        RECT 79.570 186.970 79.890 187.030 ;
        RECT 98.890 186.970 99.210 187.030 ;
        RECT 98.890 186.150 99.210 186.210 ;
        RECT 99.365 186.150 99.655 186.195 ;
        RECT 98.890 186.010 99.655 186.150 ;
        RECT 98.890 185.950 99.210 186.010 ;
        RECT 99.365 185.965 99.655 186.010 ;
      LAYER via ;
        RECT 79.600 186.970 79.860 187.230 ;
        RECT 98.920 186.970 99.180 187.230 ;
        RECT 98.920 185.950 99.180 186.210 ;
      LAYER met2 ;
        RECT 79.580 189.615 79.880 190.005 ;
        RECT 79.590 187.950 79.870 189.615 ;
        RECT 79.660 187.260 79.800 187.950 ;
        RECT 79.600 186.940 79.860 187.260 ;
        RECT 98.920 186.940 99.180 187.260 ;
        RECT 98.980 186.240 99.120 186.940 ;
        RECT 98.920 185.920 99.180 186.240 ;
      LAYER via2 ;
        RECT 79.580 189.660 79.880 189.960 ;
      LAYER met3 ;
        RECT 77.490 224.760 77.990 225.760 ;
        RECT 77.590 210.950 77.890 224.760 ;
        RECT 77.590 210.650 79.880 210.950 ;
        RECT 79.580 190.190 79.880 210.650 ;
        RECT 79.380 189.430 80.080 190.190 ;
      LAYER via3 ;
        RECT 77.540 224.810 77.940 225.710 ;
      LAYER met4 ;
        RECT 77.490 224.760 77.990 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER li1 ;
        RECT 85.155 185.875 85.415 186.335 ;
        RECT 86.015 185.875 86.275 186.335 ;
        RECT 85.155 185.705 86.275 185.875 ;
        RECT 85.155 185.455 85.415 185.705 ;
        RECT 84.660 185.285 85.415 185.455 ;
        RECT 84.660 184.775 85.065 185.285 ;
        RECT 84.660 184.605 86.310 184.775 ;
        RECT 85.155 184.215 85.415 184.605 ;
        RECT 86.015 184.215 86.310 184.605 ;
      LAYER mcon ;
        RECT 85.165 185.995 85.335 186.165 ;
      LAYER met1 ;
        RECT 77.730 186.150 78.050 186.210 ;
        RECT 85.105 186.150 85.395 186.195 ;
        RECT 77.730 186.010 85.395 186.150 ;
        RECT 77.730 185.950 78.050 186.010 ;
        RECT 85.105 185.965 85.395 186.010 ;
      LAYER via ;
        RECT 77.760 185.950 78.020 186.210 ;
      LAYER met2 ;
        RECT 77.740 189.615 78.040 190.005 ;
        RECT 77.750 187.950 78.030 189.615 ;
        RECT 77.820 186.240 77.960 187.950 ;
        RECT 77.760 185.920 78.020 186.240 ;
      LAYER via2 ;
        RECT 77.740 189.660 78.040 189.960 ;
      LAYER met3 ;
        RECT 73.810 224.760 74.310 225.760 ;
        RECT 73.910 209.950 74.210 224.760 ;
        RECT 73.910 209.650 78.040 209.950 ;
        RECT 77.740 190.190 78.040 209.650 ;
        RECT 77.540 189.430 78.240 190.190 ;
      LAYER via3 ;
        RECT 73.860 224.810 74.260 225.710 ;
      LAYER met4 ;
        RECT 73.810 224.760 74.310 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 77.265 185.430 77.520 186.335 ;
        RECT 77.265 184.700 77.435 185.430 ;
        RECT 77.265 184.125 77.520 184.700 ;
      LAYER mcon ;
        RECT 77.345 185.995 77.515 186.165 ;
      LAYER met1 ;
        RECT 75.890 186.150 76.210 186.210 ;
        RECT 77.285 186.150 77.575 186.195 ;
        RECT 75.890 186.010 77.575 186.150 ;
        RECT 75.890 185.950 76.210 186.010 ;
        RECT 77.285 185.965 77.575 186.010 ;
      LAYER via ;
        RECT 75.920 185.950 76.180 186.210 ;
      LAYER met2 ;
        RECT 75.900 189.615 76.200 190.005 ;
        RECT 75.910 187.950 76.190 189.615 ;
        RECT 75.980 186.240 76.120 187.950 ;
        RECT 75.920 185.920 76.180 186.240 ;
      LAYER via2 ;
        RECT 75.900 189.660 76.200 189.960 ;
      LAYER met3 ;
        RECT 70.130 224.760 70.630 225.760 ;
        RECT 70.230 208.950 70.530 224.760 ;
        RECT 70.230 208.650 76.200 208.950 ;
        RECT 75.900 190.190 76.200 208.650 ;
        RECT 75.700 189.430 76.400 190.190 ;
      LAYER via3 ;
        RECT 70.180 224.810 70.580 225.710 ;
      LAYER met4 ;
        RECT 70.130 224.760 70.630 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 74.965 185.430 75.220 186.335 ;
        RECT 74.965 184.700 75.135 185.430 ;
        RECT 74.965 184.125 75.220 184.700 ;
      LAYER mcon ;
        RECT 75.045 185.995 75.215 186.165 ;
      LAYER met1 ;
        RECT 74.050 186.150 74.370 186.210 ;
        RECT 74.985 186.150 75.275 186.195 ;
        RECT 74.050 186.010 75.275 186.150 ;
        RECT 74.050 185.950 74.370 186.010 ;
        RECT 74.985 185.965 75.275 186.010 ;
      LAYER via ;
        RECT 74.080 185.950 74.340 186.210 ;
      LAYER met2 ;
        RECT 74.060 189.615 74.360 190.005 ;
        RECT 74.070 187.950 74.350 189.615 ;
        RECT 74.140 186.240 74.280 187.950 ;
        RECT 74.080 185.920 74.340 186.240 ;
      LAYER via2 ;
        RECT 74.060 189.660 74.360 189.960 ;
      LAYER met3 ;
        RECT 66.450 224.760 66.950 225.760 ;
        RECT 66.550 207.950 66.850 224.760 ;
        RECT 66.550 207.650 74.360 207.950 ;
        RECT 74.060 190.190 74.360 207.650 ;
        RECT 73.860 189.430 74.560 190.190 ;
      LAYER via3 ;
        RECT 66.500 224.810 66.900 225.710 ;
      LAYER met4 ;
        RECT 66.450 224.760 66.950 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 72.205 185.430 72.460 186.335 ;
        RECT 72.205 184.700 72.375 185.430 ;
        RECT 72.205 184.125 72.460 184.700 ;
      LAYER mcon ;
        RECT 72.285 185.995 72.455 186.165 ;
      LAYER met1 ;
        RECT 72.210 185.950 72.530 186.210 ;
      LAYER via ;
        RECT 72.240 185.950 72.500 186.210 ;
      LAYER met2 ;
        RECT 72.220 189.615 72.520 190.005 ;
        RECT 72.230 187.950 72.510 189.615 ;
        RECT 72.300 186.240 72.440 187.950 ;
        RECT 72.240 185.920 72.500 186.240 ;
      LAYER via2 ;
        RECT 72.220 189.660 72.520 189.960 ;
      LAYER met3 ;
        RECT 62.770 224.760 63.270 225.760 ;
        RECT 62.870 206.950 63.170 224.760 ;
        RECT 62.870 206.650 72.520 206.950 ;
        RECT 72.220 190.190 72.520 206.650 ;
        RECT 72.020 189.430 72.720 190.190 ;
      LAYER via3 ;
        RECT 62.820 224.810 63.220 225.710 ;
      LAYER met4 ;
        RECT 62.770 224.760 63.270 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 41.590 185.175 116.030 186.780 ;
        RECT 41.590 179.735 116.030 182.565 ;
        RECT 41.590 174.295 116.030 177.125 ;
        RECT 41.590 168.855 116.030 171.685 ;
        RECT 41.590 163.415 116.030 166.245 ;
        RECT 41.590 157.975 116.030 160.805 ;
        RECT 31.560 128.360 127.040 129.790 ;
        RECT 31.560 39.010 32.990 128.360 ;
        RECT 62.250 120.980 73.910 121.790 ;
        RECT 84.910 120.980 96.570 121.790 ;
        RECT 107.570 120.980 119.230 121.790 ;
        RECT 57.650 118.730 73.910 120.980 ;
        RECT 80.310 118.730 96.570 120.980 ;
        RECT 102.970 118.730 119.230 120.980 ;
        RECT 62.250 112.010 73.910 118.730 ;
        RECT 84.910 112.010 96.570 118.730 ;
        RECT 107.570 112.010 119.230 118.730 ;
        RECT 62.250 111.030 73.930 112.010 ;
        RECT 84.910 111.030 96.590 112.010 ;
        RECT 107.570 111.030 119.250 112.010 ;
        RECT 39.590 103.640 51.250 104.450 ;
        RECT 62.250 103.640 73.910 104.450 ;
        RECT 84.910 103.640 96.570 104.450 ;
        RECT 107.570 103.640 119.230 104.450 ;
        RECT 34.990 101.390 51.250 103.640 ;
        RECT 57.650 101.390 73.910 103.640 ;
        RECT 80.310 101.390 96.570 103.640 ;
        RECT 102.970 101.390 119.230 103.640 ;
        RECT 39.590 94.670 51.250 101.390 ;
        RECT 62.250 94.670 73.910 101.390 ;
        RECT 84.910 94.670 96.570 101.390 ;
        RECT 107.570 94.670 119.230 101.390 ;
        RECT 39.590 93.690 51.270 94.670 ;
        RECT 62.250 93.690 73.930 94.670 ;
        RECT 84.910 93.690 96.590 94.670 ;
        RECT 107.570 93.690 119.250 94.670 ;
        RECT 39.590 86.300 51.250 87.110 ;
        RECT 62.250 86.300 73.910 87.110 ;
        RECT 84.910 86.300 96.570 87.110 ;
        RECT 107.570 86.300 119.230 87.110 ;
        RECT 34.990 84.050 51.250 86.300 ;
        RECT 57.650 84.050 73.910 86.300 ;
        RECT 80.310 84.050 96.570 86.300 ;
        RECT 102.970 84.050 119.230 86.300 ;
        RECT 39.590 77.330 51.250 84.050 ;
        RECT 62.250 77.330 73.910 84.050 ;
        RECT 84.910 77.330 96.570 84.050 ;
        RECT 107.570 77.330 119.230 84.050 ;
        RECT 39.590 76.350 51.270 77.330 ;
        RECT 62.250 76.350 73.930 77.330 ;
        RECT 84.910 76.350 96.590 77.330 ;
        RECT 107.570 76.350 119.250 77.330 ;
        RECT 39.590 68.960 51.250 69.770 ;
        RECT 62.250 68.960 73.910 69.770 ;
        RECT 84.910 68.960 96.570 69.770 ;
        RECT 107.570 68.960 119.230 69.770 ;
        RECT 34.990 66.710 51.250 68.960 ;
        RECT 57.650 66.710 73.910 68.960 ;
        RECT 80.310 66.710 96.570 68.960 ;
        RECT 102.970 66.710 119.230 68.960 ;
        RECT 39.590 59.990 51.250 66.710 ;
        RECT 62.250 59.990 73.910 66.710 ;
        RECT 84.910 59.990 96.570 66.710 ;
        RECT 107.570 59.990 119.230 66.710 ;
        RECT 39.590 59.010 51.270 59.990 ;
        RECT 62.250 59.010 73.930 59.990 ;
        RECT 84.910 59.010 96.590 59.990 ;
        RECT 107.570 59.010 119.250 59.990 ;
        RECT 39.590 41.990 51.250 51.770 ;
        RECT 62.250 41.990 73.910 51.770 ;
        RECT 84.910 41.990 96.570 51.770 ;
        RECT 107.570 41.990 119.230 51.770 ;
        RECT 39.590 41.010 51.270 41.990 ;
        RECT 62.250 41.010 73.930 41.990 ;
        RECT 84.910 41.010 96.590 41.990 ;
        RECT 107.570 41.010 119.250 41.990 ;
        RECT 125.610 39.010 127.040 128.360 ;
        RECT 31.560 37.580 127.040 39.010 ;
      LAYER li1 ;
        RECT 41.780 186.505 115.840 186.675 ;
        RECT 41.865 185.415 43.075 186.505 ;
        RECT 44.645 185.705 44.955 186.505 ;
        RECT 45.555 186.045 45.810 186.505 ;
        RECT 46.415 185.635 46.700 186.505 ;
        RECT 48.320 185.745 48.650 186.505 ;
        RECT 42.555 184.875 43.075 185.415 ;
        RECT 49.250 185.355 49.510 186.505 ;
        RECT 50.620 185.745 50.950 186.505 ;
        RECT 51.550 185.355 51.810 186.505 ;
        RECT 52.460 185.745 52.790 186.505 ;
        RECT 53.390 185.355 53.650 186.505 ;
        RECT 54.745 185.340 55.035 186.505 ;
        RECT 55.210 185.355 55.470 186.505 ;
        RECT 56.070 185.745 56.400 186.505 ;
        RECT 57.980 185.745 58.310 186.505 ;
        RECT 58.910 185.355 59.170 186.505 ;
        RECT 59.820 185.745 60.150 186.505 ;
        RECT 60.750 185.355 61.010 186.505 ;
        RECT 61.190 185.355 61.450 186.505 ;
        RECT 62.050 185.745 62.380 186.505 ;
        RECT 63.505 185.705 63.815 186.505 ;
        RECT 64.415 186.045 64.670 186.505 ;
        RECT 65.275 185.635 65.560 186.505 ;
        RECT 66.260 185.745 66.590 186.505 ;
        RECT 67.190 185.355 67.450 186.505 ;
        RECT 67.625 185.340 67.915 186.505 ;
        RECT 68.090 185.355 68.350 186.505 ;
        RECT 68.950 185.745 69.280 186.505 ;
        RECT 70.400 185.745 70.730 186.505 ;
        RECT 71.330 185.355 71.590 186.505 ;
        RECT 71.770 185.355 72.030 186.505 ;
        RECT 72.630 185.745 72.960 186.505 ;
        RECT 74.530 185.355 74.790 186.505 ;
        RECT 75.390 185.745 75.720 186.505 ;
        RECT 76.830 185.355 77.090 186.505 ;
        RECT 77.690 185.745 78.020 186.505 ;
        RECT 78.665 185.415 80.335 186.505 ;
        RECT 79.585 184.895 80.335 185.415 ;
        RECT 80.505 185.340 80.795 186.505 ;
        RECT 82.035 185.355 82.365 186.505 ;
        RECT 82.875 185.705 83.205 186.505 ;
        RECT 83.725 185.705 83.965 186.505 ;
        RECT 84.700 185.635 84.985 186.505 ;
        RECT 85.590 186.045 85.845 186.505 ;
        RECT 86.445 185.705 86.755 186.505 ;
        RECT 87.845 185.745 88.175 186.505 ;
        RECT 89.685 185.745 90.015 186.505 ;
        RECT 91.525 185.745 91.855 186.505 ;
        RECT 93.385 185.340 93.675 186.505 ;
        RECT 93.855 185.355 94.185 186.505 ;
        RECT 94.695 185.705 95.025 186.505 ;
        RECT 95.535 185.705 95.865 186.505 ;
        RECT 96.385 185.705 96.625 186.505 ;
        RECT 97.295 185.355 97.465 186.505 ;
        RECT 98.960 185.635 99.245 186.505 ;
        RECT 99.850 186.045 100.105 186.505 ;
        RECT 100.705 185.705 101.015 186.505 ;
        RECT 102.415 185.745 102.585 186.505 ;
        RECT 104.955 185.365 105.125 186.505 ;
        RECT 106.265 185.340 106.555 186.505 ;
        RECT 107.650 185.355 107.910 186.505 ;
        RECT 108.510 185.745 108.840 186.505 ;
        RECT 109.995 185.365 110.165 186.505 ;
        RECT 112.535 185.745 112.705 186.505 ;
        RECT 114.545 185.415 115.755 186.505 ;
        RECT 114.545 184.875 115.065 185.415 ;
        RECT 42.555 182.325 43.075 182.865 ;
        RECT 41.865 181.235 43.075 182.325 ;
        RECT 44.170 181.235 44.430 182.385 ;
        RECT 45.030 181.235 45.360 181.995 ;
        RECT 46.480 181.235 46.810 181.995 ;
        RECT 47.410 181.235 47.670 182.385 ;
        RECT 51.250 181.670 51.600 182.920 ;
        RECT 61.625 182.325 63.315 182.845 ;
        RECT 54.705 181.915 55.035 182.105 ;
        RECT 47.845 181.235 53.190 181.670 ;
        RECT 53.365 181.235 53.625 181.745 ;
        RECT 54.705 181.740 54.900 181.915 ;
        RECT 54.285 181.235 54.900 181.740 ;
        RECT 55.715 181.235 55.930 181.780 ;
        RECT 56.600 181.235 56.925 182.220 ;
        RECT 57.925 181.235 58.775 181.685 ;
        RECT 59.375 181.235 59.630 182.235 ;
        RECT 59.805 181.235 63.315 182.325 ;
        RECT 64.235 181.235 64.405 181.995 ;
        RECT 66.775 181.235 66.945 182.375 ;
        RECT 67.625 181.235 67.915 182.400 ;
        RECT 69.755 181.235 69.925 181.995 ;
        RECT 72.295 181.235 72.465 182.375 ;
        RECT 73.895 181.235 74.065 181.995 ;
        RECT 76.435 181.235 76.605 182.375 ;
        RECT 77.715 181.235 78.100 181.660 ;
        RECT 79.130 181.235 79.515 181.660 ;
        RECT 80.725 181.235 81.110 181.660 ;
        RECT 82.395 181.235 82.565 182.375 ;
        RECT 86.945 182.325 87.695 182.845 ;
        RECT 84.935 181.235 85.105 181.995 ;
        RECT 86.025 181.235 87.695 182.325 ;
        RECT 88.375 181.235 88.545 182.375 ;
        RECT 90.915 181.235 91.085 181.995 ;
        RECT 92.445 181.235 92.775 181.995 ;
        RECT 93.385 181.235 93.675 182.400 ;
        RECT 94.355 181.235 94.525 182.375 ;
        RECT 96.895 181.235 97.065 181.995 ;
        RECT 98.495 181.235 98.665 182.375 ;
        RECT 101.035 181.235 101.205 181.995 ;
        RECT 102.595 181.235 102.925 182.385 ;
        RECT 103.435 181.235 103.765 182.035 ;
        RECT 104.275 181.235 104.605 182.035 ;
        RECT 105.125 181.235 105.365 182.035 ;
        RECT 106.035 181.235 106.205 182.385 ;
        RECT 107.235 181.235 107.405 182.375 ;
        RECT 109.775 181.235 109.945 181.995 ;
        RECT 111.375 181.235 111.615 182.035 ;
        RECT 112.135 181.235 112.465 182.035 ;
        RECT 112.975 181.235 113.305 182.385 ;
        RECT 114.545 182.325 115.065 182.865 ;
        RECT 114.545 181.235 115.755 182.325 ;
        RECT 41.780 181.065 115.840 181.235 ;
        RECT 41.865 179.975 43.075 181.065 ;
        RECT 43.245 180.630 48.590 181.065 ;
        RECT 50.195 180.635 50.605 181.065 ;
        RECT 51.350 180.645 51.680 181.065 ;
        RECT 42.555 179.435 43.075 179.975 ;
        RECT 46.650 179.380 47.000 180.630 ;
        RECT 52.650 179.965 52.980 181.065 ;
        RECT 53.425 179.925 53.635 181.065 ;
        RECT 54.305 179.925 54.535 181.065 ;
        RECT 54.745 179.900 55.035 181.065 ;
        RECT 55.205 180.630 60.550 181.065 ;
        RECT 58.610 179.380 58.960 180.630 ;
        RECT 60.725 179.975 62.395 181.065 ;
        RECT 61.645 179.455 62.395 179.975 ;
        RECT 63.535 179.925 63.705 181.065 ;
        RECT 66.075 180.305 66.245 181.065 ;
        RECT 68.525 180.305 68.855 181.065 ;
        RECT 69.465 179.975 70.675 181.065 ;
        RECT 70.945 180.605 71.155 181.065 ;
        RECT 71.825 180.265 71.995 181.065 ;
        RECT 70.155 179.435 70.675 179.975 ;
        RECT 72.665 179.925 72.930 181.065 ;
        RECT 73.145 179.975 74.815 181.065 ;
        RECT 74.990 180.640 75.325 181.065 ;
        RECT 75.885 180.285 76.215 181.065 ;
        RECT 76.825 179.975 80.335 181.065 ;
        RECT 74.065 179.455 74.815 179.975 ;
        RECT 78.645 179.455 80.335 179.975 ;
        RECT 80.505 179.900 80.795 181.065 ;
        RECT 80.965 180.630 86.310 181.065 ;
        RECT 84.370 179.380 84.720 180.630 ;
        RECT 86.485 179.975 88.155 181.065 ;
        RECT 89.535 180.305 89.705 181.065 ;
        RECT 87.405 179.455 88.155 179.975 ;
        RECT 92.075 179.925 92.245 181.065 ;
        RECT 93.365 180.305 93.695 181.065 ;
        RECT 95.230 179.915 95.490 181.065 ;
        RECT 96.090 180.305 96.420 181.065 ;
        RECT 97.505 180.305 97.835 181.065 ;
        RECT 98.885 180.305 99.215 181.065 ;
        RECT 100.795 179.925 100.965 181.065 ;
        RECT 103.335 180.305 103.505 181.065 ;
        RECT 104.865 180.305 105.195 181.065 ;
        RECT 106.265 179.900 106.555 181.065 ;
        RECT 107.165 180.285 107.495 181.065 ;
        RECT 108.055 180.640 108.390 181.065 ;
        RECT 109.630 180.640 110.015 181.065 ;
        RECT 111.225 180.640 111.610 181.065 ;
        RECT 112.640 180.640 113.025 181.065 ;
        RECT 114.545 179.975 115.755 181.065 ;
        RECT 114.545 179.435 115.065 179.975 ;
        RECT 42.555 176.885 43.075 177.425 ;
        RECT 41.865 175.795 43.075 176.885 ;
        RECT 46.650 176.230 47.000 177.480 ;
        RECT 43.245 175.795 48.590 176.230 ;
        RECT 50.135 175.795 50.845 176.570 ;
        RECT 51.935 175.795 52.265 176.515 ;
        RECT 55.850 176.230 56.200 177.480 ;
        RECT 52.445 175.795 57.790 176.230 ;
        RECT 58.935 175.795 59.105 176.935 ;
        RECT 66.245 176.885 66.995 177.405 ;
        RECT 61.475 175.795 61.645 176.555 ;
        RECT 63.045 175.795 63.355 176.595 ;
        RECT 63.955 175.795 64.210 176.255 ;
        RECT 64.815 175.795 65.100 176.665 ;
        RECT 65.325 175.795 66.995 176.885 ;
        RECT 67.625 175.795 67.915 176.960 ;
        RECT 68.190 175.795 68.445 176.595 ;
        RECT 69.115 175.795 69.285 176.595 ;
        RECT 69.955 175.795 70.215 176.935 ;
        RECT 73.790 176.230 74.140 177.480 ;
        RECT 70.385 175.795 75.730 176.230 ;
        RECT 76.415 175.795 76.585 176.935 ;
        RECT 92.695 176.885 93.215 177.425 ;
        RECT 78.955 175.795 79.125 176.555 ;
        RECT 80.475 175.795 80.805 176.175 ;
        RECT 83.290 175.795 83.640 176.175 ;
        RECT 84.230 175.795 84.560 176.175 ;
        RECT 86.055 175.795 86.385 176.175 ;
        RECT 88.775 175.795 89.105 176.175 ;
        RECT 90.355 175.795 90.685 176.515 ;
        RECT 91.355 175.795 91.635 176.465 ;
        RECT 92.005 175.795 93.215 176.885 ;
        RECT 93.385 175.795 93.675 176.960 ;
        RECT 94.355 175.795 94.525 176.935 ;
        RECT 96.895 175.795 97.065 176.555 ;
        RECT 98.335 175.795 98.505 176.945 ;
        RECT 99.175 175.795 99.415 176.595 ;
        RECT 99.935 175.795 100.265 176.595 ;
        RECT 100.775 175.795 101.105 176.595 ;
        RECT 101.615 175.795 101.945 176.945 ;
        RECT 103.555 175.795 103.725 176.935 ;
        RECT 106.095 175.795 106.265 176.555 ;
        RECT 107.650 175.795 107.910 176.945 ;
        RECT 108.510 175.795 108.840 176.555 ;
        RECT 110.415 175.795 110.745 176.945 ;
        RECT 111.255 175.795 111.585 176.595 ;
        RECT 112.095 175.795 112.425 176.595 ;
        RECT 112.945 175.795 113.185 176.595 ;
        RECT 113.855 175.795 114.025 176.945 ;
        RECT 114.545 176.885 115.065 177.425 ;
        RECT 114.545 175.795 115.755 176.885 ;
        RECT 41.780 175.625 115.840 175.795 ;
        RECT 41.865 174.535 43.075 175.625 ;
        RECT 43.245 175.190 48.590 175.625 ;
        RECT 42.555 173.995 43.075 174.535 ;
        RECT 46.650 173.940 47.000 175.190 ;
        RECT 48.765 175.115 49.065 175.625 ;
        RECT 49.735 175.115 50.365 175.625 ;
        RECT 51.495 175.115 51.795 175.625 ;
        RECT 51.985 174.535 54.575 175.625 ;
        RECT 53.365 174.015 54.575 174.535 ;
        RECT 54.745 174.460 55.035 175.625 ;
        RECT 55.205 175.115 55.505 175.625 ;
        RECT 56.175 175.115 56.805 175.625 ;
        RECT 57.935 175.115 58.235 175.625 ;
        RECT 59.075 174.905 59.405 175.625 ;
        RECT 60.075 174.955 60.355 175.625 ;
        RECT 60.725 174.535 61.935 175.625 ;
        RECT 62.855 174.865 63.025 175.625 ;
        RECT 61.415 173.995 61.935 174.535 ;
        RECT 65.395 174.485 65.565 175.625 ;
        RECT 66.755 174.485 66.925 175.625 ;
        RECT 69.295 174.865 69.465 175.625 ;
        RECT 70.815 175.245 71.145 175.625 ;
        RECT 73.535 175.245 73.865 175.625 ;
        RECT 75.360 175.245 75.690 175.625 ;
        RECT 76.280 175.245 76.630 175.625 ;
        RECT 79.115 175.245 79.445 175.625 ;
        RECT 80.505 174.460 80.795 175.625 ;
        RECT 81.715 174.865 81.885 175.625 ;
        RECT 84.255 174.485 84.425 175.625 ;
        RECT 85.545 174.865 85.875 175.625 ;
        RECT 86.485 174.535 88.155 175.625 ;
        RECT 89.075 174.865 89.245 175.625 ;
        RECT 87.405 174.015 88.155 174.535 ;
        RECT 91.615 174.485 91.785 175.625 ;
        RECT 93.215 174.865 93.385 175.625 ;
        RECT 95.755 174.485 95.925 175.625 ;
        RECT 98.035 174.485 98.205 175.625 ;
        RECT 100.575 174.865 100.745 175.625 ;
        RECT 102.175 174.485 102.345 175.625 ;
        RECT 104.715 174.865 104.885 175.625 ;
        RECT 106.265 174.460 106.555 175.625 ;
        RECT 107.235 174.485 107.405 175.625 ;
        RECT 109.775 174.865 109.945 175.625 ;
        RECT 111.935 174.475 112.265 175.625 ;
        RECT 112.775 174.825 113.105 175.625 ;
        RECT 113.625 174.825 113.865 175.625 ;
        RECT 114.545 174.535 115.755 175.625 ;
        RECT 114.545 173.995 115.065 174.535 ;
        RECT 42.555 171.445 43.075 171.985 ;
        RECT 41.865 170.355 43.075 171.445 ;
        RECT 46.650 170.790 47.000 172.040 ;
        RECT 52.170 170.790 52.520 172.040 ;
        RECT 55.205 171.445 55.955 171.965 ;
        RECT 43.245 170.355 48.590 170.790 ;
        RECT 48.765 170.355 54.110 170.790 ;
        RECT 54.285 170.355 55.955 171.445 ;
        RECT 56.635 170.355 56.805 171.495 ;
        RECT 61.185 171.445 61.935 171.965 ;
        RECT 66.935 171.445 67.455 171.985 ;
        RECT 59.175 170.355 59.345 171.115 ;
        RECT 60.265 170.355 61.935 171.445 ;
        RECT 63.435 170.355 63.685 171.275 ;
        RECT 65.035 170.355 65.365 171.145 ;
        RECT 66.245 170.355 67.455 171.445 ;
        RECT 67.625 170.355 67.915 171.520 ;
        RECT 68.525 170.355 68.855 171.115 ;
        RECT 72.870 170.790 73.220 172.040 ;
        RECT 78.390 170.790 78.740 172.040 ;
        RECT 69.465 170.355 74.810 170.790 ;
        RECT 74.985 170.355 80.330 170.790 ;
        RECT 81.475 170.355 81.645 171.495 ;
        RECT 84.015 170.355 84.185 171.115 ;
        RECT 87.060 170.355 87.390 170.735 ;
        RECT 88.785 170.355 89.115 171.535 ;
        RECT 92.005 171.445 92.755 171.965 ;
        RECT 89.815 170.355 89.985 171.195 ;
        RECT 90.655 170.355 90.865 171.195 ;
        RECT 91.085 170.355 92.755 171.445 ;
        RECT 93.385 170.355 93.675 171.520 ;
        RECT 95.225 171.445 96.435 171.965 ;
        RECT 93.845 170.355 96.435 171.445 ;
        RECT 98.100 170.355 98.430 170.735 ;
        RECT 99.825 170.355 100.155 171.535 ;
        RECT 103.505 171.445 104.715 171.965 ;
        RECT 100.855 170.355 101.025 171.195 ;
        RECT 101.695 170.355 101.905 171.195 ;
        RECT 102.125 170.355 104.715 171.445 ;
        RECT 114.545 171.445 115.065 171.985 ;
        RECT 105.315 170.355 105.645 170.735 ;
        RECT 108.035 170.355 108.365 170.735 ;
        RECT 109.860 170.355 110.190 170.735 ;
        RECT 110.780 170.355 111.130 170.735 ;
        RECT 113.615 170.355 113.945 170.735 ;
        RECT 114.545 170.355 115.755 171.445 ;
        RECT 41.780 170.185 115.840 170.355 ;
        RECT 41.865 169.095 43.075 170.185 ;
        RECT 43.245 169.750 48.590 170.185 ;
        RECT 48.765 169.750 54.110 170.185 ;
        RECT 42.555 168.555 43.075 169.095 ;
        RECT 46.650 168.500 47.000 169.750 ;
        RECT 52.170 168.500 52.520 169.750 ;
        RECT 54.745 169.020 55.035 170.185 ;
        RECT 55.205 169.095 58.715 170.185 ;
        RECT 58.885 169.095 60.095 170.185 ;
        RECT 61.015 169.425 61.185 170.185 ;
        RECT 57.025 168.575 58.715 169.095 ;
        RECT 59.575 168.555 60.095 169.095 ;
        RECT 63.555 169.045 63.725 170.185 ;
        RECT 64.405 169.095 66.995 170.185 ;
        RECT 68.515 169.725 68.845 170.185 ;
        RECT 70.075 169.385 70.400 170.185 ;
        RECT 65.785 168.575 66.995 169.095 ;
        RECT 71.325 169.045 71.595 170.185 ;
        RECT 72.275 169.045 72.445 170.185 ;
        RECT 74.815 169.425 74.985 170.185 ;
        RECT 75.905 169.095 79.415 170.185 ;
        RECT 77.725 168.575 79.415 169.095 ;
        RECT 80.505 169.020 80.795 170.185 ;
        RECT 82.315 169.805 82.645 170.185 ;
        RECT 85.035 169.805 85.365 170.185 ;
        RECT 86.860 169.805 87.190 170.185 ;
        RECT 87.780 169.805 88.130 170.185 ;
        RECT 90.615 169.805 90.945 170.185 ;
        RECT 93.355 169.725 93.685 170.185 ;
        RECT 94.915 169.385 95.240 170.185 ;
        RECT 96.165 169.045 96.435 170.185 ;
        RECT 97.035 169.805 97.365 170.185 ;
        RECT 99.755 169.805 100.085 170.185 ;
        RECT 101.580 169.805 101.910 170.185 ;
        RECT 102.500 169.805 102.850 170.185 ;
        RECT 105.335 169.805 105.665 170.185 ;
        RECT 106.265 169.020 106.555 170.185 ;
        RECT 107.235 169.045 107.405 170.185 ;
        RECT 109.775 169.425 109.945 170.185 ;
        RECT 111.305 169.425 111.635 170.185 ;
        RECT 112.685 169.425 113.015 170.185 ;
        RECT 114.545 169.095 115.755 170.185 ;
        RECT 114.545 168.555 115.065 169.095 ;
        RECT 42.555 166.005 43.075 166.545 ;
        RECT 41.865 164.915 43.075 166.005 ;
        RECT 46.650 165.350 47.000 166.600 ;
        RECT 49.685 166.005 50.435 166.525 ;
        RECT 43.245 164.915 48.590 165.350 ;
        RECT 48.765 164.915 50.435 166.005 ;
        RECT 63.670 165.350 64.020 166.600 ;
        RECT 66.705 166.005 67.455 166.525 ;
        RECT 51.035 164.915 51.365 165.295 ;
        RECT 53.850 164.915 54.200 165.295 ;
        RECT 54.790 164.915 55.120 165.295 ;
        RECT 56.615 164.915 56.945 165.295 ;
        RECT 59.335 164.915 59.665 165.295 ;
        RECT 60.265 164.915 65.610 165.350 ;
        RECT 65.785 164.915 67.455 166.005 ;
        RECT 67.625 164.915 67.915 166.080 ;
        RECT 69.465 166.005 70.675 166.525 ;
        RECT 73.605 166.005 74.355 166.525 ;
        RECT 78.895 166.005 79.415 166.545 ;
        RECT 68.085 164.915 70.675 166.005 ;
        RECT 70.850 164.915 71.185 165.340 ;
        RECT 71.745 164.915 72.075 165.695 ;
        RECT 72.685 164.915 74.355 166.005 ;
        RECT 75.395 164.915 75.645 165.835 ;
        RECT 76.995 164.915 77.325 165.705 ;
        RECT 78.205 164.915 79.415 166.005 ;
        RECT 79.590 164.915 79.925 165.340 ;
        RECT 80.485 164.915 80.815 165.695 ;
        RECT 84.830 165.350 85.180 166.600 ;
        RECT 88.765 166.005 90.455 166.525 ;
        RECT 81.425 164.915 86.770 165.350 ;
        RECT 86.945 164.915 90.455 166.005 ;
        RECT 91.550 164.915 91.885 165.340 ;
        RECT 92.445 164.915 92.775 165.695 ;
        RECT 93.385 164.915 93.675 166.080 ;
        RECT 94.735 164.915 95.065 165.375 ;
        RECT 96.295 164.915 96.620 165.715 ;
        RECT 97.545 164.915 97.815 166.055 ;
        RECT 101.390 165.350 101.740 166.600 ;
        RECT 97.985 164.915 103.330 165.350 ;
        RECT 104.475 164.915 104.685 165.755 ;
        RECT 105.355 164.915 105.525 165.755 ;
        RECT 106.225 164.915 106.555 166.095 ;
        RECT 107.950 164.915 108.280 165.295 ;
        RECT 110.455 164.915 110.625 166.055 ;
        RECT 114.545 166.005 115.065 166.545 ;
        RECT 112.995 164.915 113.165 165.675 ;
        RECT 114.545 164.915 115.755 166.005 ;
        RECT 41.780 164.745 115.840 164.915 ;
        RECT 41.865 163.655 43.075 164.745 ;
        RECT 43.245 164.310 48.590 164.745 ;
        RECT 48.765 164.310 54.110 164.745 ;
        RECT 42.555 163.115 43.075 163.655 ;
        RECT 46.650 163.060 47.000 164.310 ;
        RECT 52.170 163.060 52.520 164.310 ;
        RECT 54.745 163.580 55.035 164.745 ;
        RECT 55.225 164.235 55.525 164.745 ;
        RECT 56.655 164.235 57.285 164.745 ;
        RECT 57.955 164.235 58.255 164.745 ;
        RECT 58.425 163.655 61.015 164.745 ;
        RECT 61.615 164.365 61.945 164.745 ;
        RECT 64.430 164.365 64.780 164.745 ;
        RECT 65.370 164.365 65.700 164.745 ;
        RECT 67.195 164.365 67.525 164.745 ;
        RECT 69.915 164.365 70.245 164.745 ;
        RECT 70.845 164.310 76.190 164.745 ;
        RECT 59.805 163.135 61.015 163.655 ;
        RECT 74.250 163.060 74.600 164.310 ;
        RECT 76.365 163.655 78.035 164.745 ;
        RECT 78.670 164.320 79.005 164.745 ;
        RECT 79.565 163.965 79.895 164.745 ;
        RECT 77.285 163.135 78.035 163.655 ;
        RECT 80.505 163.580 80.795 164.745 ;
        RECT 81.855 164.285 82.185 164.745 ;
        RECT 83.415 163.945 83.740 164.745 ;
        RECT 84.665 163.605 84.935 164.745 ;
        RECT 86.535 163.605 86.705 164.745 ;
        RECT 89.075 163.985 89.245 164.745 ;
        RECT 90.165 163.655 93.675 164.745 ;
        RECT 91.985 163.135 93.675 163.655 ;
        RECT 94.355 163.605 94.525 164.745 ;
        RECT 96.895 163.985 97.065 164.745 ;
        RECT 98.495 163.605 98.665 164.745 ;
        RECT 101.035 163.985 101.205 164.745 ;
        RECT 102.565 163.965 102.895 164.745 ;
        RECT 103.455 164.320 103.790 164.745 ;
        RECT 103.965 163.655 105.635 164.745 ;
        RECT 104.885 163.135 105.635 163.655 ;
        RECT 106.265 163.580 106.555 164.745 ;
        RECT 106.725 163.655 109.315 164.745 ;
        RECT 109.925 163.985 110.255 164.745 ;
        RECT 111.305 163.985 111.635 164.745 ;
        RECT 112.685 163.985 113.015 164.745 ;
        RECT 108.105 163.135 109.315 163.655 ;
        RECT 114.545 163.655 115.755 164.745 ;
        RECT 114.545 163.115 115.065 163.655 ;
        RECT 42.555 160.565 43.075 161.105 ;
        RECT 41.865 159.475 43.075 160.565 ;
        RECT 46.650 159.910 47.000 161.160 ;
        RECT 50.145 160.565 51.355 161.085 ;
        RECT 59.805 160.565 61.015 161.085 ;
        RECT 43.245 159.475 48.590 159.910 ;
        RECT 48.765 159.475 51.355 160.565 ;
        RECT 52.955 159.475 53.125 160.325 ;
        RECT 53.795 159.475 53.965 159.985 ;
        RECT 55.205 159.475 55.505 159.985 ;
        RECT 56.175 159.475 56.805 159.985 ;
        RECT 57.935 159.475 58.235 159.985 ;
        RECT 58.425 159.475 61.015 160.565 ;
        RECT 61.185 159.475 61.485 159.985 ;
        RECT 62.155 159.475 62.785 159.985 ;
        RECT 63.915 159.475 64.215 159.985 ;
        RECT 65.375 159.475 65.545 160.325 ;
        RECT 66.215 159.475 66.385 159.985 ;
        RECT 67.625 159.475 67.915 160.640 ;
        RECT 69.005 160.565 69.755 161.085 ;
        RECT 68.085 159.475 69.755 160.565 ;
        RECT 70.435 159.475 70.605 160.615 ;
        RECT 72.975 159.475 73.145 160.235 ;
        RECT 74.575 159.475 74.745 160.615 ;
        RECT 77.115 159.475 77.285 160.235 ;
        RECT 79.125 159.475 79.425 159.985 ;
        RECT 80.095 159.475 80.725 159.985 ;
        RECT 81.855 159.475 82.155 159.985 ;
        RECT 85.750 159.910 86.100 161.160 ;
        RECT 88.785 160.565 89.535 161.085 ;
        RECT 82.345 159.475 87.690 159.910 ;
        RECT 87.865 159.475 89.535 160.565 ;
        RECT 90.775 159.475 90.945 159.985 ;
        RECT 91.615 159.475 91.785 160.325 ;
        RECT 93.385 159.475 93.675 160.640 ;
        RECT 94.765 160.565 95.515 161.085 ;
        RECT 99.345 160.565 101.035 161.085 ;
        RECT 93.845 159.475 95.515 160.565 ;
        RECT 95.690 159.475 96.025 159.900 ;
        RECT 96.585 159.475 96.915 160.255 ;
        RECT 97.525 159.475 101.035 160.565 ;
        RECT 102.175 159.475 102.345 160.615 ;
        RECT 110.175 160.565 110.695 161.105 ;
        RECT 104.715 159.475 104.885 160.235 ;
        RECT 106.515 159.475 106.845 160.265 ;
        RECT 108.195 159.475 108.445 160.395 ;
        RECT 109.485 159.475 110.695 160.565 ;
        RECT 114.545 160.565 115.065 161.105 ;
        RECT 111.305 159.475 111.635 160.235 ;
        RECT 112.685 159.475 113.015 160.235 ;
        RECT 114.545 159.475 115.755 160.565 ;
        RECT 41.780 159.305 115.840 159.475 ;
        RECT 41.865 158.215 43.075 159.305 ;
        RECT 44.145 158.545 44.475 159.305 ;
        RECT 45.085 158.215 48.595 159.305 ;
        RECT 49.205 158.545 49.535 159.305 ;
        RECT 50.145 158.215 53.655 159.305 ;
        RECT 42.555 157.675 43.075 158.215 ;
        RECT 46.905 157.695 48.595 158.215 ;
        RECT 51.965 157.695 53.655 158.215 ;
        RECT 54.745 158.140 55.035 159.305 ;
        RECT 55.645 158.545 55.975 159.305 ;
        RECT 56.585 158.215 58.255 159.305 ;
        RECT 59.325 158.545 59.655 159.305 ;
        RECT 60.265 158.215 63.775 159.305 ;
        RECT 64.385 158.545 64.715 159.305 ;
        RECT 65.325 158.215 66.995 159.305 ;
        RECT 57.505 157.695 58.255 158.215 ;
        RECT 62.085 157.695 63.775 158.215 ;
        RECT 66.245 157.695 66.995 158.215 ;
        RECT 67.625 158.140 67.915 159.305 ;
        RECT 68.085 158.795 68.385 159.305 ;
        RECT 69.055 158.795 69.685 159.305 ;
        RECT 70.815 158.795 71.115 159.305 ;
        RECT 71.745 158.545 72.075 159.305 ;
        RECT 72.685 158.215 73.895 159.305 ;
        RECT 74.505 158.545 74.835 159.305 ;
        RECT 75.445 158.215 78.955 159.305 ;
        RECT 79.565 158.545 79.895 159.305 ;
        RECT 73.375 157.675 73.895 158.215 ;
        RECT 77.265 157.695 78.955 158.215 ;
        RECT 80.505 158.140 80.795 159.305 ;
        RECT 80.965 158.215 82.635 159.305 ;
        RECT 83.285 158.795 83.585 159.305 ;
        RECT 84.715 158.795 85.345 159.305 ;
        RECT 86.015 158.795 86.315 159.305 ;
        RECT 86.925 158.545 87.255 159.305 ;
        RECT 87.865 158.215 89.075 159.305 ;
        RECT 89.685 158.545 90.015 159.305 ;
        RECT 90.625 158.215 93.215 159.305 ;
        RECT 81.885 157.695 82.635 158.215 ;
        RECT 88.555 157.675 89.075 158.215 ;
        RECT 92.005 157.695 93.215 158.215 ;
        RECT 93.385 158.140 93.675 159.305 ;
        RECT 94.745 158.545 95.075 159.305 ;
        RECT 95.685 158.215 99.195 159.305 ;
        RECT 99.805 158.545 100.135 159.305 ;
        RECT 100.745 158.215 104.255 159.305 ;
        RECT 104.865 158.545 105.195 159.305 ;
        RECT 97.505 157.695 99.195 158.215 ;
        RECT 102.565 157.695 104.255 158.215 ;
        RECT 106.265 158.140 106.555 159.305 ;
        RECT 107.615 158.845 107.945 159.305 ;
        RECT 109.175 158.505 109.500 159.305 ;
        RECT 110.425 158.165 110.695 159.305 ;
        RECT 111.305 158.545 111.635 159.305 ;
        RECT 113.605 158.545 113.935 159.305 ;
        RECT 114.545 158.215 115.755 159.305 ;
        RECT 114.545 157.675 115.065 158.215 ;
        RECT 31.845 129.335 126.755 129.505 ;
        RECT 31.845 38.035 32.015 129.335 ;
        RECT 59.470 119.460 59.640 120.500 ;
        RECT 60.870 119.460 61.040 120.500 ;
        RECT 58.040 119.060 58.410 119.270 ;
        RECT 67.700 117.270 67.870 121.310 ;
        RECT 68.290 117.270 68.460 121.310 ;
        RECT 70.170 117.270 70.340 121.310 ;
        RECT 72.050 117.270 72.220 121.310 ;
        RECT 76.540 119.360 76.890 121.520 ;
        RECT 82.130 119.460 82.300 120.500 ;
        RECT 83.530 119.460 83.700 120.500 ;
        RECT 80.700 119.060 81.070 119.270 ;
        RECT 90.360 117.270 90.530 121.310 ;
        RECT 90.950 117.270 91.120 121.310 ;
        RECT 92.830 117.270 93.000 121.310 ;
        RECT 94.710 117.270 94.880 121.310 ;
        RECT 99.200 119.360 99.550 121.520 ;
        RECT 104.790 119.460 104.960 120.500 ;
        RECT 106.190 119.460 106.360 120.500 ;
        RECT 103.360 119.060 103.730 119.270 ;
        RECT 113.020 117.270 113.190 121.310 ;
        RECT 113.610 117.270 113.780 121.310 ;
        RECT 115.490 117.270 115.660 121.310 ;
        RECT 117.370 117.270 117.540 121.310 ;
        RECT 121.860 119.360 122.210 121.520 ;
        RECT 67.700 112.090 67.870 116.130 ;
        RECT 68.290 112.090 68.460 116.130 ;
        RECT 70.170 112.090 70.340 116.130 ;
        RECT 72.050 112.090 72.220 116.130 ;
        RECT 90.360 112.090 90.530 116.130 ;
        RECT 90.950 112.090 91.120 116.130 ;
        RECT 92.830 112.090 93.000 116.130 ;
        RECT 94.710 112.090 94.880 116.130 ;
        RECT 113.020 112.090 113.190 116.130 ;
        RECT 113.610 112.090 113.780 116.130 ;
        RECT 115.490 112.090 115.660 116.130 ;
        RECT 117.370 112.090 117.540 116.130 ;
        RECT 64.190 111.400 64.400 111.770 ;
        RECT 66.070 111.400 66.280 111.770 ;
        RECT 67.950 111.400 68.160 111.770 ;
        RECT 69.830 111.400 70.040 111.770 ;
        RECT 71.710 111.400 71.920 111.770 ;
        RECT 86.850 111.400 87.060 111.770 ;
        RECT 88.730 111.400 88.940 111.770 ;
        RECT 90.610 111.400 90.820 111.770 ;
        RECT 92.490 111.400 92.700 111.770 ;
        RECT 94.370 111.400 94.580 111.770 ;
        RECT 109.510 111.400 109.720 111.770 ;
        RECT 111.390 111.400 111.600 111.770 ;
        RECT 113.270 111.400 113.480 111.770 ;
        RECT 115.150 111.400 115.360 111.770 ;
        RECT 117.030 111.400 117.240 111.770 ;
        RECT 56.220 107.280 56.570 109.440 ;
        RECT 36.810 102.120 36.980 103.160 ;
        RECT 38.210 102.120 38.380 103.160 ;
        RECT 35.380 101.720 35.750 101.930 ;
        RECT 45.040 99.930 45.210 103.970 ;
        RECT 45.630 99.930 45.800 103.970 ;
        RECT 47.510 99.930 47.680 103.970 ;
        RECT 49.390 99.930 49.560 103.970 ;
        RECT 53.880 102.020 54.230 104.180 ;
        RECT 59.470 102.120 59.640 103.160 ;
        RECT 60.870 102.120 61.040 103.160 ;
        RECT 58.040 101.720 58.410 101.930 ;
        RECT 67.700 99.930 67.870 103.970 ;
        RECT 68.290 99.930 68.460 103.970 ;
        RECT 70.170 99.930 70.340 103.970 ;
        RECT 72.050 99.930 72.220 103.970 ;
        RECT 76.540 102.020 76.890 104.180 ;
        RECT 82.130 102.120 82.300 103.160 ;
        RECT 83.530 102.120 83.700 103.160 ;
        RECT 80.700 101.720 81.070 101.930 ;
        RECT 90.360 99.930 90.530 103.970 ;
        RECT 90.950 99.930 91.120 103.970 ;
        RECT 92.830 99.930 93.000 103.970 ;
        RECT 94.710 99.930 94.880 103.970 ;
        RECT 99.200 102.020 99.550 104.180 ;
        RECT 104.790 102.120 104.960 103.160 ;
        RECT 106.190 102.120 106.360 103.160 ;
        RECT 103.360 101.720 103.730 101.930 ;
        RECT 113.020 99.930 113.190 103.970 ;
        RECT 113.610 99.930 113.780 103.970 ;
        RECT 115.490 99.930 115.660 103.970 ;
        RECT 117.370 99.930 117.540 103.970 ;
        RECT 121.860 102.020 122.210 104.180 ;
        RECT 45.040 94.750 45.210 98.790 ;
        RECT 45.630 94.750 45.800 98.790 ;
        RECT 47.510 94.750 47.680 98.790 ;
        RECT 49.390 94.750 49.560 98.790 ;
        RECT 67.700 94.750 67.870 98.790 ;
        RECT 68.290 94.750 68.460 98.790 ;
        RECT 70.170 94.750 70.340 98.790 ;
        RECT 72.050 94.750 72.220 98.790 ;
        RECT 90.360 94.750 90.530 98.790 ;
        RECT 90.950 94.750 91.120 98.790 ;
        RECT 92.830 94.750 93.000 98.790 ;
        RECT 94.710 94.750 94.880 98.790 ;
        RECT 113.020 94.750 113.190 98.790 ;
        RECT 113.610 94.750 113.780 98.790 ;
        RECT 115.490 94.750 115.660 98.790 ;
        RECT 117.370 94.750 117.540 98.790 ;
        RECT 41.530 94.060 41.740 94.430 ;
        RECT 43.410 94.060 43.620 94.430 ;
        RECT 45.290 94.060 45.500 94.430 ;
        RECT 47.170 94.060 47.380 94.430 ;
        RECT 49.050 94.060 49.260 94.430 ;
        RECT 64.190 94.060 64.400 94.430 ;
        RECT 66.070 94.060 66.280 94.430 ;
        RECT 67.950 94.060 68.160 94.430 ;
        RECT 69.830 94.060 70.040 94.430 ;
        RECT 71.710 94.060 71.920 94.430 ;
        RECT 86.850 94.060 87.060 94.430 ;
        RECT 88.730 94.060 88.940 94.430 ;
        RECT 90.610 94.060 90.820 94.430 ;
        RECT 92.490 94.060 92.700 94.430 ;
        RECT 94.370 94.060 94.580 94.430 ;
        RECT 109.510 94.060 109.720 94.430 ;
        RECT 111.390 94.060 111.600 94.430 ;
        RECT 113.270 94.060 113.480 94.430 ;
        RECT 115.150 94.060 115.360 94.430 ;
        RECT 117.030 94.060 117.240 94.430 ;
        RECT 36.810 84.780 36.980 85.820 ;
        RECT 38.210 84.780 38.380 85.820 ;
        RECT 35.380 84.380 35.750 84.590 ;
        RECT 45.040 82.590 45.210 86.630 ;
        RECT 45.630 82.590 45.800 86.630 ;
        RECT 47.510 82.590 47.680 86.630 ;
        RECT 49.390 82.590 49.560 86.630 ;
        RECT 53.880 84.680 54.230 86.840 ;
        RECT 59.470 84.780 59.640 85.820 ;
        RECT 60.870 84.780 61.040 85.820 ;
        RECT 58.040 84.380 58.410 84.590 ;
        RECT 67.700 82.590 67.870 86.630 ;
        RECT 68.290 82.590 68.460 86.630 ;
        RECT 70.170 82.590 70.340 86.630 ;
        RECT 72.050 82.590 72.220 86.630 ;
        RECT 76.540 84.680 76.890 86.840 ;
        RECT 82.130 84.780 82.300 85.820 ;
        RECT 83.530 84.780 83.700 85.820 ;
        RECT 80.700 84.380 81.070 84.590 ;
        RECT 90.360 82.590 90.530 86.630 ;
        RECT 90.950 82.590 91.120 86.630 ;
        RECT 92.830 82.590 93.000 86.630 ;
        RECT 94.710 82.590 94.880 86.630 ;
        RECT 99.200 84.680 99.550 86.840 ;
        RECT 104.790 84.780 104.960 85.820 ;
        RECT 106.190 84.780 106.360 85.820 ;
        RECT 103.360 84.380 103.730 84.590 ;
        RECT 113.020 82.590 113.190 86.630 ;
        RECT 113.610 82.590 113.780 86.630 ;
        RECT 115.490 82.590 115.660 86.630 ;
        RECT 117.370 82.590 117.540 86.630 ;
        RECT 121.860 84.680 122.210 86.840 ;
        RECT 45.040 77.410 45.210 81.450 ;
        RECT 45.630 77.410 45.800 81.450 ;
        RECT 47.510 77.410 47.680 81.450 ;
        RECT 49.390 77.410 49.560 81.450 ;
        RECT 67.700 77.410 67.870 81.450 ;
        RECT 68.290 77.410 68.460 81.450 ;
        RECT 70.170 77.410 70.340 81.450 ;
        RECT 72.050 77.410 72.220 81.450 ;
        RECT 90.360 77.410 90.530 81.450 ;
        RECT 90.950 77.410 91.120 81.450 ;
        RECT 92.830 77.410 93.000 81.450 ;
        RECT 94.710 77.410 94.880 81.450 ;
        RECT 113.020 77.410 113.190 81.450 ;
        RECT 113.610 77.410 113.780 81.450 ;
        RECT 115.490 77.410 115.660 81.450 ;
        RECT 117.370 77.410 117.540 81.450 ;
        RECT 41.530 76.720 41.740 77.090 ;
        RECT 43.410 76.720 43.620 77.090 ;
        RECT 45.290 76.720 45.500 77.090 ;
        RECT 47.170 76.720 47.380 77.090 ;
        RECT 49.050 76.720 49.260 77.090 ;
        RECT 64.190 76.720 64.400 77.090 ;
        RECT 66.070 76.720 66.280 77.090 ;
        RECT 67.950 76.720 68.160 77.090 ;
        RECT 69.830 76.720 70.040 77.090 ;
        RECT 71.710 76.720 71.920 77.090 ;
        RECT 86.850 76.720 87.060 77.090 ;
        RECT 88.730 76.720 88.940 77.090 ;
        RECT 90.610 76.720 90.820 77.090 ;
        RECT 92.490 76.720 92.700 77.090 ;
        RECT 94.370 76.720 94.580 77.090 ;
        RECT 109.510 76.720 109.720 77.090 ;
        RECT 111.390 76.720 111.600 77.090 ;
        RECT 113.270 76.720 113.480 77.090 ;
        RECT 115.150 76.720 115.360 77.090 ;
        RECT 117.030 76.720 117.240 77.090 ;
        RECT 36.810 67.440 36.980 68.480 ;
        RECT 38.210 67.440 38.380 68.480 ;
        RECT 35.380 67.040 35.750 67.250 ;
        RECT 45.040 65.250 45.210 69.290 ;
        RECT 45.630 65.250 45.800 69.290 ;
        RECT 47.510 65.250 47.680 69.290 ;
        RECT 49.390 65.250 49.560 69.290 ;
        RECT 53.880 67.340 54.230 69.500 ;
        RECT 59.470 67.440 59.640 68.480 ;
        RECT 60.870 67.440 61.040 68.480 ;
        RECT 58.040 67.040 58.410 67.250 ;
        RECT 67.700 65.250 67.870 69.290 ;
        RECT 68.290 65.250 68.460 69.290 ;
        RECT 70.170 65.250 70.340 69.290 ;
        RECT 72.050 65.250 72.220 69.290 ;
        RECT 76.540 67.340 76.890 69.500 ;
        RECT 82.130 67.440 82.300 68.480 ;
        RECT 83.530 67.440 83.700 68.480 ;
        RECT 80.700 67.040 81.070 67.250 ;
        RECT 90.360 65.250 90.530 69.290 ;
        RECT 90.950 65.250 91.120 69.290 ;
        RECT 92.830 65.250 93.000 69.290 ;
        RECT 94.710 65.250 94.880 69.290 ;
        RECT 99.200 67.340 99.550 69.500 ;
        RECT 104.790 67.440 104.960 68.480 ;
        RECT 106.190 67.440 106.360 68.480 ;
        RECT 103.360 67.040 103.730 67.250 ;
        RECT 113.020 65.250 113.190 69.290 ;
        RECT 113.610 65.250 113.780 69.290 ;
        RECT 115.490 65.250 115.660 69.290 ;
        RECT 117.370 65.250 117.540 69.290 ;
        RECT 121.860 67.340 122.210 69.500 ;
        RECT 45.040 60.070 45.210 64.110 ;
        RECT 45.630 60.070 45.800 64.110 ;
        RECT 47.510 60.070 47.680 64.110 ;
        RECT 49.390 60.070 49.560 64.110 ;
        RECT 67.700 60.070 67.870 64.110 ;
        RECT 68.290 60.070 68.460 64.110 ;
        RECT 70.170 60.070 70.340 64.110 ;
        RECT 72.050 60.070 72.220 64.110 ;
        RECT 90.360 60.070 90.530 64.110 ;
        RECT 90.950 60.070 91.120 64.110 ;
        RECT 92.830 60.070 93.000 64.110 ;
        RECT 94.710 60.070 94.880 64.110 ;
        RECT 113.020 60.070 113.190 64.110 ;
        RECT 113.610 60.070 113.780 64.110 ;
        RECT 115.490 60.070 115.660 64.110 ;
        RECT 117.370 60.070 117.540 64.110 ;
        RECT 41.530 59.380 41.740 59.750 ;
        RECT 43.410 59.380 43.620 59.750 ;
        RECT 45.290 59.380 45.500 59.750 ;
        RECT 47.170 59.380 47.380 59.750 ;
        RECT 49.050 59.380 49.260 59.750 ;
        RECT 64.190 59.380 64.400 59.750 ;
        RECT 66.070 59.380 66.280 59.750 ;
        RECT 67.950 59.380 68.160 59.750 ;
        RECT 69.830 59.380 70.040 59.750 ;
        RECT 71.710 59.380 71.920 59.750 ;
        RECT 86.850 59.380 87.060 59.750 ;
        RECT 88.730 59.380 88.940 59.750 ;
        RECT 90.610 59.380 90.820 59.750 ;
        RECT 92.490 59.380 92.700 59.750 ;
        RECT 94.370 59.380 94.580 59.750 ;
        RECT 109.510 59.380 109.720 59.750 ;
        RECT 111.390 59.380 111.600 59.750 ;
        RECT 113.270 59.380 113.480 59.750 ;
        RECT 115.150 59.380 115.360 59.750 ;
        RECT 117.030 59.380 117.240 59.750 ;
        RECT 45.040 47.250 45.210 51.290 ;
        RECT 45.630 47.250 45.800 51.290 ;
        RECT 47.510 47.250 47.680 51.290 ;
        RECT 49.390 47.250 49.560 51.290 ;
        RECT 53.880 49.340 54.230 51.500 ;
        RECT 67.700 47.250 67.870 51.290 ;
        RECT 68.290 47.250 68.460 51.290 ;
        RECT 70.170 47.250 70.340 51.290 ;
        RECT 72.050 47.250 72.220 51.290 ;
        RECT 76.540 49.340 76.890 51.500 ;
        RECT 90.360 47.250 90.530 51.290 ;
        RECT 90.950 47.250 91.120 51.290 ;
        RECT 92.830 47.250 93.000 51.290 ;
        RECT 94.710 47.250 94.880 51.290 ;
        RECT 99.200 49.340 99.550 51.500 ;
        RECT 113.020 47.250 113.190 51.290 ;
        RECT 113.610 47.250 113.780 51.290 ;
        RECT 115.490 47.250 115.660 51.290 ;
        RECT 117.370 47.250 117.540 51.290 ;
        RECT 121.860 49.340 122.210 51.500 ;
        RECT 45.040 42.070 45.210 46.110 ;
        RECT 45.630 42.070 45.800 46.110 ;
        RECT 47.510 42.070 47.680 46.110 ;
        RECT 49.390 42.070 49.560 46.110 ;
        RECT 67.700 42.070 67.870 46.110 ;
        RECT 68.290 42.070 68.460 46.110 ;
        RECT 70.170 42.070 70.340 46.110 ;
        RECT 72.050 42.070 72.220 46.110 ;
        RECT 90.360 42.070 90.530 46.110 ;
        RECT 90.950 42.070 91.120 46.110 ;
        RECT 92.830 42.070 93.000 46.110 ;
        RECT 94.710 42.070 94.880 46.110 ;
        RECT 113.020 42.070 113.190 46.110 ;
        RECT 113.610 42.070 113.780 46.110 ;
        RECT 115.490 42.070 115.660 46.110 ;
        RECT 117.370 42.070 117.540 46.110 ;
        RECT 41.530 41.380 41.740 41.750 ;
        RECT 43.410 41.380 43.620 41.750 ;
        RECT 45.290 41.380 45.500 41.750 ;
        RECT 47.170 41.380 47.380 41.750 ;
        RECT 49.050 41.380 49.260 41.750 ;
        RECT 64.190 41.380 64.400 41.750 ;
        RECT 66.070 41.380 66.280 41.750 ;
        RECT 67.950 41.380 68.160 41.750 ;
        RECT 69.830 41.380 70.040 41.750 ;
        RECT 71.710 41.380 71.920 41.750 ;
        RECT 86.850 41.380 87.060 41.750 ;
        RECT 88.730 41.380 88.940 41.750 ;
        RECT 90.610 41.380 90.820 41.750 ;
        RECT 92.490 41.380 92.700 41.750 ;
        RECT 94.370 41.380 94.580 41.750 ;
        RECT 109.510 41.380 109.720 41.750 ;
        RECT 111.390 41.380 111.600 41.750 ;
        RECT 113.270 41.380 113.480 41.750 ;
        RECT 115.150 41.380 115.360 41.750 ;
        RECT 117.030 41.380 117.240 41.750 ;
        RECT 126.585 38.035 126.755 129.335 ;
        RECT 31.845 37.865 126.755 38.035 ;
      LAYER mcon ;
        RECT 41.925 186.505 42.095 186.675 ;
        RECT 42.385 186.505 42.555 186.675 ;
        RECT 42.845 186.505 43.015 186.675 ;
        RECT 43.305 186.505 43.475 186.675 ;
        RECT 43.765 186.505 43.935 186.675 ;
        RECT 44.225 186.505 44.395 186.675 ;
        RECT 44.685 186.505 44.855 186.675 ;
        RECT 45.145 186.505 45.315 186.675 ;
        RECT 45.605 186.505 45.775 186.675 ;
        RECT 46.065 186.505 46.235 186.675 ;
        RECT 46.525 186.505 46.695 186.675 ;
        RECT 46.985 186.505 47.155 186.675 ;
        RECT 47.445 186.505 47.615 186.675 ;
        RECT 47.905 186.505 48.075 186.675 ;
        RECT 48.365 186.505 48.535 186.675 ;
        RECT 48.825 186.505 48.995 186.675 ;
        RECT 49.285 186.505 49.455 186.675 ;
        RECT 49.745 186.505 49.915 186.675 ;
        RECT 50.205 186.505 50.375 186.675 ;
        RECT 50.665 186.505 50.835 186.675 ;
        RECT 51.125 186.505 51.295 186.675 ;
        RECT 51.585 186.505 51.755 186.675 ;
        RECT 52.045 186.505 52.215 186.675 ;
        RECT 52.505 186.505 52.675 186.675 ;
        RECT 52.965 186.505 53.135 186.675 ;
        RECT 53.425 186.505 53.595 186.675 ;
        RECT 53.885 186.505 54.055 186.675 ;
        RECT 54.345 186.505 54.515 186.675 ;
        RECT 54.805 186.505 54.975 186.675 ;
        RECT 55.265 186.505 55.435 186.675 ;
        RECT 55.725 186.505 55.895 186.675 ;
        RECT 56.185 186.505 56.355 186.675 ;
        RECT 56.645 186.505 56.815 186.675 ;
        RECT 57.105 186.505 57.275 186.675 ;
        RECT 57.565 186.505 57.735 186.675 ;
        RECT 58.025 186.505 58.195 186.675 ;
        RECT 58.485 186.505 58.655 186.675 ;
        RECT 58.945 186.505 59.115 186.675 ;
        RECT 59.405 186.505 59.575 186.675 ;
        RECT 59.865 186.505 60.035 186.675 ;
        RECT 60.325 186.505 60.495 186.675 ;
        RECT 60.785 186.505 60.955 186.675 ;
        RECT 61.245 186.505 61.415 186.675 ;
        RECT 61.705 186.505 61.875 186.675 ;
        RECT 62.165 186.505 62.335 186.675 ;
        RECT 62.625 186.505 62.795 186.675 ;
        RECT 63.085 186.505 63.255 186.675 ;
        RECT 63.545 186.505 63.715 186.675 ;
        RECT 64.005 186.505 64.175 186.675 ;
        RECT 64.465 186.505 64.635 186.675 ;
        RECT 64.925 186.505 65.095 186.675 ;
        RECT 65.385 186.505 65.555 186.675 ;
        RECT 65.845 186.505 66.015 186.675 ;
        RECT 66.305 186.505 66.475 186.675 ;
        RECT 66.765 186.505 66.935 186.675 ;
        RECT 67.225 186.505 67.395 186.675 ;
        RECT 67.685 186.505 67.855 186.675 ;
        RECT 68.145 186.505 68.315 186.675 ;
        RECT 68.605 186.505 68.775 186.675 ;
        RECT 69.065 186.505 69.235 186.675 ;
        RECT 69.525 186.505 69.695 186.675 ;
        RECT 69.985 186.505 70.155 186.675 ;
        RECT 70.445 186.505 70.615 186.675 ;
        RECT 70.905 186.505 71.075 186.675 ;
        RECT 71.365 186.505 71.535 186.675 ;
        RECT 71.825 186.505 71.995 186.675 ;
        RECT 72.285 186.505 72.455 186.675 ;
        RECT 72.745 186.505 72.915 186.675 ;
        RECT 73.205 186.505 73.375 186.675 ;
        RECT 73.665 186.505 73.835 186.675 ;
        RECT 74.125 186.505 74.295 186.675 ;
        RECT 74.585 186.505 74.755 186.675 ;
        RECT 75.045 186.505 75.215 186.675 ;
        RECT 75.505 186.505 75.675 186.675 ;
        RECT 75.965 186.505 76.135 186.675 ;
        RECT 76.425 186.505 76.595 186.675 ;
        RECT 76.885 186.505 77.055 186.675 ;
        RECT 77.345 186.505 77.515 186.675 ;
        RECT 77.805 186.505 77.975 186.675 ;
        RECT 78.265 186.505 78.435 186.675 ;
        RECT 78.725 186.505 78.895 186.675 ;
        RECT 79.185 186.505 79.355 186.675 ;
        RECT 79.645 186.505 79.815 186.675 ;
        RECT 80.105 186.505 80.275 186.675 ;
        RECT 80.565 186.505 80.735 186.675 ;
        RECT 81.025 186.505 81.195 186.675 ;
        RECT 81.485 186.505 81.655 186.675 ;
        RECT 81.945 186.505 82.115 186.675 ;
        RECT 82.405 186.505 82.575 186.675 ;
        RECT 82.865 186.505 83.035 186.675 ;
        RECT 83.325 186.505 83.495 186.675 ;
        RECT 83.785 186.505 83.955 186.675 ;
        RECT 84.245 186.505 84.415 186.675 ;
        RECT 84.705 186.505 84.875 186.675 ;
        RECT 85.165 186.505 85.335 186.675 ;
        RECT 85.625 186.505 85.795 186.675 ;
        RECT 86.085 186.505 86.255 186.675 ;
        RECT 86.545 186.505 86.715 186.675 ;
        RECT 87.005 186.505 87.175 186.675 ;
        RECT 87.465 186.505 87.635 186.675 ;
        RECT 87.925 186.505 88.095 186.675 ;
        RECT 88.385 186.505 88.555 186.675 ;
        RECT 88.845 186.505 89.015 186.675 ;
        RECT 89.305 186.505 89.475 186.675 ;
        RECT 89.765 186.505 89.935 186.675 ;
        RECT 90.225 186.505 90.395 186.675 ;
        RECT 90.685 186.505 90.855 186.675 ;
        RECT 91.145 186.505 91.315 186.675 ;
        RECT 91.605 186.505 91.775 186.675 ;
        RECT 92.065 186.505 92.235 186.675 ;
        RECT 92.525 186.505 92.695 186.675 ;
        RECT 92.985 186.505 93.155 186.675 ;
        RECT 93.445 186.505 93.615 186.675 ;
        RECT 93.905 186.505 94.075 186.675 ;
        RECT 94.365 186.505 94.535 186.675 ;
        RECT 94.825 186.505 94.995 186.675 ;
        RECT 95.285 186.505 95.455 186.675 ;
        RECT 95.745 186.505 95.915 186.675 ;
        RECT 96.205 186.505 96.375 186.675 ;
        RECT 96.665 186.505 96.835 186.675 ;
        RECT 97.125 186.505 97.295 186.675 ;
        RECT 97.585 186.505 97.755 186.675 ;
        RECT 98.045 186.505 98.215 186.675 ;
        RECT 98.505 186.505 98.675 186.675 ;
        RECT 98.965 186.505 99.135 186.675 ;
        RECT 99.425 186.505 99.595 186.675 ;
        RECT 99.885 186.505 100.055 186.675 ;
        RECT 100.345 186.505 100.515 186.675 ;
        RECT 100.805 186.505 100.975 186.675 ;
        RECT 101.265 186.505 101.435 186.675 ;
        RECT 101.725 186.505 101.895 186.675 ;
        RECT 102.185 186.505 102.355 186.675 ;
        RECT 102.645 186.505 102.815 186.675 ;
        RECT 103.105 186.505 103.275 186.675 ;
        RECT 103.565 186.505 103.735 186.675 ;
        RECT 104.025 186.505 104.195 186.675 ;
        RECT 104.485 186.505 104.655 186.675 ;
        RECT 104.945 186.505 105.115 186.675 ;
        RECT 105.405 186.505 105.575 186.675 ;
        RECT 105.865 186.505 106.035 186.675 ;
        RECT 106.325 186.505 106.495 186.675 ;
        RECT 106.785 186.505 106.955 186.675 ;
        RECT 107.245 186.505 107.415 186.675 ;
        RECT 107.705 186.505 107.875 186.675 ;
        RECT 108.165 186.505 108.335 186.675 ;
        RECT 108.625 186.505 108.795 186.675 ;
        RECT 109.085 186.505 109.255 186.675 ;
        RECT 109.545 186.505 109.715 186.675 ;
        RECT 110.005 186.505 110.175 186.675 ;
        RECT 110.465 186.505 110.635 186.675 ;
        RECT 110.925 186.505 111.095 186.675 ;
        RECT 111.385 186.505 111.555 186.675 ;
        RECT 111.845 186.505 112.015 186.675 ;
        RECT 112.305 186.505 112.475 186.675 ;
        RECT 112.765 186.505 112.935 186.675 ;
        RECT 113.225 186.505 113.395 186.675 ;
        RECT 113.685 186.505 113.855 186.675 ;
        RECT 114.145 186.505 114.315 186.675 ;
        RECT 114.605 186.505 114.775 186.675 ;
        RECT 115.065 186.505 115.235 186.675 ;
        RECT 115.525 186.505 115.695 186.675 ;
        RECT 41.925 181.065 42.095 181.235 ;
        RECT 42.385 181.065 42.555 181.235 ;
        RECT 42.845 181.065 43.015 181.235 ;
        RECT 43.305 181.065 43.475 181.235 ;
        RECT 43.765 181.065 43.935 181.235 ;
        RECT 44.225 181.065 44.395 181.235 ;
        RECT 44.685 181.065 44.855 181.235 ;
        RECT 45.145 181.065 45.315 181.235 ;
        RECT 45.605 181.065 45.775 181.235 ;
        RECT 46.065 181.065 46.235 181.235 ;
        RECT 46.525 181.065 46.695 181.235 ;
        RECT 46.985 181.065 47.155 181.235 ;
        RECT 47.445 181.065 47.615 181.235 ;
        RECT 47.905 181.065 48.075 181.235 ;
        RECT 48.365 181.065 48.535 181.235 ;
        RECT 48.825 181.065 48.995 181.235 ;
        RECT 49.285 181.065 49.455 181.235 ;
        RECT 49.745 181.065 49.915 181.235 ;
        RECT 50.205 181.065 50.375 181.235 ;
        RECT 50.665 181.065 50.835 181.235 ;
        RECT 51.125 181.065 51.295 181.235 ;
        RECT 51.585 181.065 51.755 181.235 ;
        RECT 52.045 181.065 52.215 181.235 ;
        RECT 52.505 181.065 52.675 181.235 ;
        RECT 52.965 181.065 53.135 181.235 ;
        RECT 53.425 181.065 53.595 181.235 ;
        RECT 53.885 181.065 54.055 181.235 ;
        RECT 54.345 181.065 54.515 181.235 ;
        RECT 54.805 181.065 54.975 181.235 ;
        RECT 55.265 181.065 55.435 181.235 ;
        RECT 55.725 181.065 55.895 181.235 ;
        RECT 56.185 181.065 56.355 181.235 ;
        RECT 56.645 181.065 56.815 181.235 ;
        RECT 57.105 181.065 57.275 181.235 ;
        RECT 57.565 181.065 57.735 181.235 ;
        RECT 58.025 181.065 58.195 181.235 ;
        RECT 58.485 181.065 58.655 181.235 ;
        RECT 58.945 181.065 59.115 181.235 ;
        RECT 59.405 181.065 59.575 181.235 ;
        RECT 59.865 181.065 60.035 181.235 ;
        RECT 60.325 181.065 60.495 181.235 ;
        RECT 60.785 181.065 60.955 181.235 ;
        RECT 61.245 181.065 61.415 181.235 ;
        RECT 61.705 181.065 61.875 181.235 ;
        RECT 62.165 181.065 62.335 181.235 ;
        RECT 62.625 181.065 62.795 181.235 ;
        RECT 63.085 181.065 63.255 181.235 ;
        RECT 63.545 181.065 63.715 181.235 ;
        RECT 64.005 181.065 64.175 181.235 ;
        RECT 64.465 181.065 64.635 181.235 ;
        RECT 64.925 181.065 65.095 181.235 ;
        RECT 65.385 181.065 65.555 181.235 ;
        RECT 65.845 181.065 66.015 181.235 ;
        RECT 66.305 181.065 66.475 181.235 ;
        RECT 66.765 181.065 66.935 181.235 ;
        RECT 67.225 181.065 67.395 181.235 ;
        RECT 67.685 181.065 67.855 181.235 ;
        RECT 68.145 181.065 68.315 181.235 ;
        RECT 68.605 181.065 68.775 181.235 ;
        RECT 69.065 181.065 69.235 181.235 ;
        RECT 69.525 181.065 69.695 181.235 ;
        RECT 69.985 181.065 70.155 181.235 ;
        RECT 70.445 181.065 70.615 181.235 ;
        RECT 70.905 181.065 71.075 181.235 ;
        RECT 71.365 181.065 71.535 181.235 ;
        RECT 71.825 181.065 71.995 181.235 ;
        RECT 72.285 181.065 72.455 181.235 ;
        RECT 72.745 181.065 72.915 181.235 ;
        RECT 73.205 181.065 73.375 181.235 ;
        RECT 73.665 181.065 73.835 181.235 ;
        RECT 74.125 181.065 74.295 181.235 ;
        RECT 74.585 181.065 74.755 181.235 ;
        RECT 75.045 181.065 75.215 181.235 ;
        RECT 75.505 181.065 75.675 181.235 ;
        RECT 75.965 181.065 76.135 181.235 ;
        RECT 76.425 181.065 76.595 181.235 ;
        RECT 76.885 181.065 77.055 181.235 ;
        RECT 77.345 181.065 77.515 181.235 ;
        RECT 77.805 181.065 77.975 181.235 ;
        RECT 78.265 181.065 78.435 181.235 ;
        RECT 78.725 181.065 78.895 181.235 ;
        RECT 79.185 181.065 79.355 181.235 ;
        RECT 79.645 181.065 79.815 181.235 ;
        RECT 80.105 181.065 80.275 181.235 ;
        RECT 80.565 181.065 80.735 181.235 ;
        RECT 81.025 181.065 81.195 181.235 ;
        RECT 81.485 181.065 81.655 181.235 ;
        RECT 81.945 181.065 82.115 181.235 ;
        RECT 82.405 181.065 82.575 181.235 ;
        RECT 82.865 181.065 83.035 181.235 ;
        RECT 83.325 181.065 83.495 181.235 ;
        RECT 83.785 181.065 83.955 181.235 ;
        RECT 84.245 181.065 84.415 181.235 ;
        RECT 84.705 181.065 84.875 181.235 ;
        RECT 85.165 181.065 85.335 181.235 ;
        RECT 85.625 181.065 85.795 181.235 ;
        RECT 86.085 181.065 86.255 181.235 ;
        RECT 86.545 181.065 86.715 181.235 ;
        RECT 87.005 181.065 87.175 181.235 ;
        RECT 87.465 181.065 87.635 181.235 ;
        RECT 87.925 181.065 88.095 181.235 ;
        RECT 88.385 181.065 88.555 181.235 ;
        RECT 88.845 181.065 89.015 181.235 ;
        RECT 89.305 181.065 89.475 181.235 ;
        RECT 89.765 181.065 89.935 181.235 ;
        RECT 90.225 181.065 90.395 181.235 ;
        RECT 90.685 181.065 90.855 181.235 ;
        RECT 91.145 181.065 91.315 181.235 ;
        RECT 91.605 181.065 91.775 181.235 ;
        RECT 92.065 181.065 92.235 181.235 ;
        RECT 92.525 181.065 92.695 181.235 ;
        RECT 92.985 181.065 93.155 181.235 ;
        RECT 93.445 181.065 93.615 181.235 ;
        RECT 93.905 181.065 94.075 181.235 ;
        RECT 94.365 181.065 94.535 181.235 ;
        RECT 94.825 181.065 94.995 181.235 ;
        RECT 95.285 181.065 95.455 181.235 ;
        RECT 95.745 181.065 95.915 181.235 ;
        RECT 96.205 181.065 96.375 181.235 ;
        RECT 96.665 181.065 96.835 181.235 ;
        RECT 97.125 181.065 97.295 181.235 ;
        RECT 97.585 181.065 97.755 181.235 ;
        RECT 98.045 181.065 98.215 181.235 ;
        RECT 98.505 181.065 98.675 181.235 ;
        RECT 98.965 181.065 99.135 181.235 ;
        RECT 99.425 181.065 99.595 181.235 ;
        RECT 99.885 181.065 100.055 181.235 ;
        RECT 100.345 181.065 100.515 181.235 ;
        RECT 100.805 181.065 100.975 181.235 ;
        RECT 101.265 181.065 101.435 181.235 ;
        RECT 101.725 181.065 101.895 181.235 ;
        RECT 102.185 181.065 102.355 181.235 ;
        RECT 102.645 181.065 102.815 181.235 ;
        RECT 103.105 181.065 103.275 181.235 ;
        RECT 103.565 181.065 103.735 181.235 ;
        RECT 104.025 181.065 104.195 181.235 ;
        RECT 104.485 181.065 104.655 181.235 ;
        RECT 104.945 181.065 105.115 181.235 ;
        RECT 105.405 181.065 105.575 181.235 ;
        RECT 105.865 181.065 106.035 181.235 ;
        RECT 106.325 181.065 106.495 181.235 ;
        RECT 106.785 181.065 106.955 181.235 ;
        RECT 107.245 181.065 107.415 181.235 ;
        RECT 107.705 181.065 107.875 181.235 ;
        RECT 108.165 181.065 108.335 181.235 ;
        RECT 108.625 181.065 108.795 181.235 ;
        RECT 109.085 181.065 109.255 181.235 ;
        RECT 109.545 181.065 109.715 181.235 ;
        RECT 110.005 181.065 110.175 181.235 ;
        RECT 110.465 181.065 110.635 181.235 ;
        RECT 110.925 181.065 111.095 181.235 ;
        RECT 111.385 181.065 111.555 181.235 ;
        RECT 111.845 181.065 112.015 181.235 ;
        RECT 112.305 181.065 112.475 181.235 ;
        RECT 112.765 181.065 112.935 181.235 ;
        RECT 113.225 181.065 113.395 181.235 ;
        RECT 113.685 181.065 113.855 181.235 ;
        RECT 114.145 181.065 114.315 181.235 ;
        RECT 114.605 181.065 114.775 181.235 ;
        RECT 115.065 181.065 115.235 181.235 ;
        RECT 115.525 181.065 115.695 181.235 ;
        RECT 41.925 175.625 42.095 175.795 ;
        RECT 42.385 175.625 42.555 175.795 ;
        RECT 42.845 175.625 43.015 175.795 ;
        RECT 43.305 175.625 43.475 175.795 ;
        RECT 43.765 175.625 43.935 175.795 ;
        RECT 44.225 175.625 44.395 175.795 ;
        RECT 44.685 175.625 44.855 175.795 ;
        RECT 45.145 175.625 45.315 175.795 ;
        RECT 45.605 175.625 45.775 175.795 ;
        RECT 46.065 175.625 46.235 175.795 ;
        RECT 46.525 175.625 46.695 175.795 ;
        RECT 46.985 175.625 47.155 175.795 ;
        RECT 47.445 175.625 47.615 175.795 ;
        RECT 47.905 175.625 48.075 175.795 ;
        RECT 48.365 175.625 48.535 175.795 ;
        RECT 48.825 175.625 48.995 175.795 ;
        RECT 49.285 175.625 49.455 175.795 ;
        RECT 49.745 175.625 49.915 175.795 ;
        RECT 50.205 175.625 50.375 175.795 ;
        RECT 50.665 175.625 50.835 175.795 ;
        RECT 51.125 175.625 51.295 175.795 ;
        RECT 51.585 175.625 51.755 175.795 ;
        RECT 52.045 175.625 52.215 175.795 ;
        RECT 52.505 175.625 52.675 175.795 ;
        RECT 52.965 175.625 53.135 175.795 ;
        RECT 53.425 175.625 53.595 175.795 ;
        RECT 53.885 175.625 54.055 175.795 ;
        RECT 54.345 175.625 54.515 175.795 ;
        RECT 54.805 175.625 54.975 175.795 ;
        RECT 55.265 175.625 55.435 175.795 ;
        RECT 55.725 175.625 55.895 175.795 ;
        RECT 56.185 175.625 56.355 175.795 ;
        RECT 56.645 175.625 56.815 175.795 ;
        RECT 57.105 175.625 57.275 175.795 ;
        RECT 57.565 175.625 57.735 175.795 ;
        RECT 58.025 175.625 58.195 175.795 ;
        RECT 58.485 175.625 58.655 175.795 ;
        RECT 58.945 175.625 59.115 175.795 ;
        RECT 59.405 175.625 59.575 175.795 ;
        RECT 59.865 175.625 60.035 175.795 ;
        RECT 60.325 175.625 60.495 175.795 ;
        RECT 60.785 175.625 60.955 175.795 ;
        RECT 61.245 175.625 61.415 175.795 ;
        RECT 61.705 175.625 61.875 175.795 ;
        RECT 62.165 175.625 62.335 175.795 ;
        RECT 62.625 175.625 62.795 175.795 ;
        RECT 63.085 175.625 63.255 175.795 ;
        RECT 63.545 175.625 63.715 175.795 ;
        RECT 64.005 175.625 64.175 175.795 ;
        RECT 64.465 175.625 64.635 175.795 ;
        RECT 64.925 175.625 65.095 175.795 ;
        RECT 65.385 175.625 65.555 175.795 ;
        RECT 65.845 175.625 66.015 175.795 ;
        RECT 66.305 175.625 66.475 175.795 ;
        RECT 66.765 175.625 66.935 175.795 ;
        RECT 67.225 175.625 67.395 175.795 ;
        RECT 67.685 175.625 67.855 175.795 ;
        RECT 68.145 175.625 68.315 175.795 ;
        RECT 68.605 175.625 68.775 175.795 ;
        RECT 69.065 175.625 69.235 175.795 ;
        RECT 69.525 175.625 69.695 175.795 ;
        RECT 69.985 175.625 70.155 175.795 ;
        RECT 70.445 175.625 70.615 175.795 ;
        RECT 70.905 175.625 71.075 175.795 ;
        RECT 71.365 175.625 71.535 175.795 ;
        RECT 71.825 175.625 71.995 175.795 ;
        RECT 72.285 175.625 72.455 175.795 ;
        RECT 72.745 175.625 72.915 175.795 ;
        RECT 73.205 175.625 73.375 175.795 ;
        RECT 73.665 175.625 73.835 175.795 ;
        RECT 74.125 175.625 74.295 175.795 ;
        RECT 74.585 175.625 74.755 175.795 ;
        RECT 75.045 175.625 75.215 175.795 ;
        RECT 75.505 175.625 75.675 175.795 ;
        RECT 75.965 175.625 76.135 175.795 ;
        RECT 76.425 175.625 76.595 175.795 ;
        RECT 76.885 175.625 77.055 175.795 ;
        RECT 77.345 175.625 77.515 175.795 ;
        RECT 77.805 175.625 77.975 175.795 ;
        RECT 78.265 175.625 78.435 175.795 ;
        RECT 78.725 175.625 78.895 175.795 ;
        RECT 79.185 175.625 79.355 175.795 ;
        RECT 79.645 175.625 79.815 175.795 ;
        RECT 80.105 175.625 80.275 175.795 ;
        RECT 80.565 175.625 80.735 175.795 ;
        RECT 81.025 175.625 81.195 175.795 ;
        RECT 81.485 175.625 81.655 175.795 ;
        RECT 81.945 175.625 82.115 175.795 ;
        RECT 82.405 175.625 82.575 175.795 ;
        RECT 82.865 175.625 83.035 175.795 ;
        RECT 83.325 175.625 83.495 175.795 ;
        RECT 83.785 175.625 83.955 175.795 ;
        RECT 84.245 175.625 84.415 175.795 ;
        RECT 84.705 175.625 84.875 175.795 ;
        RECT 85.165 175.625 85.335 175.795 ;
        RECT 85.625 175.625 85.795 175.795 ;
        RECT 86.085 175.625 86.255 175.795 ;
        RECT 86.545 175.625 86.715 175.795 ;
        RECT 87.005 175.625 87.175 175.795 ;
        RECT 87.465 175.625 87.635 175.795 ;
        RECT 87.925 175.625 88.095 175.795 ;
        RECT 88.385 175.625 88.555 175.795 ;
        RECT 88.845 175.625 89.015 175.795 ;
        RECT 89.305 175.625 89.475 175.795 ;
        RECT 89.765 175.625 89.935 175.795 ;
        RECT 90.225 175.625 90.395 175.795 ;
        RECT 90.685 175.625 90.855 175.795 ;
        RECT 91.145 175.625 91.315 175.795 ;
        RECT 91.605 175.625 91.775 175.795 ;
        RECT 92.065 175.625 92.235 175.795 ;
        RECT 92.525 175.625 92.695 175.795 ;
        RECT 92.985 175.625 93.155 175.795 ;
        RECT 93.445 175.625 93.615 175.795 ;
        RECT 93.905 175.625 94.075 175.795 ;
        RECT 94.365 175.625 94.535 175.795 ;
        RECT 94.825 175.625 94.995 175.795 ;
        RECT 95.285 175.625 95.455 175.795 ;
        RECT 95.745 175.625 95.915 175.795 ;
        RECT 96.205 175.625 96.375 175.795 ;
        RECT 96.665 175.625 96.835 175.795 ;
        RECT 97.125 175.625 97.295 175.795 ;
        RECT 97.585 175.625 97.755 175.795 ;
        RECT 98.045 175.625 98.215 175.795 ;
        RECT 98.505 175.625 98.675 175.795 ;
        RECT 98.965 175.625 99.135 175.795 ;
        RECT 99.425 175.625 99.595 175.795 ;
        RECT 99.885 175.625 100.055 175.795 ;
        RECT 100.345 175.625 100.515 175.795 ;
        RECT 100.805 175.625 100.975 175.795 ;
        RECT 101.265 175.625 101.435 175.795 ;
        RECT 101.725 175.625 101.895 175.795 ;
        RECT 102.185 175.625 102.355 175.795 ;
        RECT 102.645 175.625 102.815 175.795 ;
        RECT 103.105 175.625 103.275 175.795 ;
        RECT 103.565 175.625 103.735 175.795 ;
        RECT 104.025 175.625 104.195 175.795 ;
        RECT 104.485 175.625 104.655 175.795 ;
        RECT 104.945 175.625 105.115 175.795 ;
        RECT 105.405 175.625 105.575 175.795 ;
        RECT 105.865 175.625 106.035 175.795 ;
        RECT 106.325 175.625 106.495 175.795 ;
        RECT 106.785 175.625 106.955 175.795 ;
        RECT 107.245 175.625 107.415 175.795 ;
        RECT 107.705 175.625 107.875 175.795 ;
        RECT 108.165 175.625 108.335 175.795 ;
        RECT 108.625 175.625 108.795 175.795 ;
        RECT 109.085 175.625 109.255 175.795 ;
        RECT 109.545 175.625 109.715 175.795 ;
        RECT 110.005 175.625 110.175 175.795 ;
        RECT 110.465 175.625 110.635 175.795 ;
        RECT 110.925 175.625 111.095 175.795 ;
        RECT 111.385 175.625 111.555 175.795 ;
        RECT 111.845 175.625 112.015 175.795 ;
        RECT 112.305 175.625 112.475 175.795 ;
        RECT 112.765 175.625 112.935 175.795 ;
        RECT 113.225 175.625 113.395 175.795 ;
        RECT 113.685 175.625 113.855 175.795 ;
        RECT 114.145 175.625 114.315 175.795 ;
        RECT 114.605 175.625 114.775 175.795 ;
        RECT 115.065 175.625 115.235 175.795 ;
        RECT 115.525 175.625 115.695 175.795 ;
        RECT 41.925 170.185 42.095 170.355 ;
        RECT 42.385 170.185 42.555 170.355 ;
        RECT 42.845 170.185 43.015 170.355 ;
        RECT 43.305 170.185 43.475 170.355 ;
        RECT 43.765 170.185 43.935 170.355 ;
        RECT 44.225 170.185 44.395 170.355 ;
        RECT 44.685 170.185 44.855 170.355 ;
        RECT 45.145 170.185 45.315 170.355 ;
        RECT 45.605 170.185 45.775 170.355 ;
        RECT 46.065 170.185 46.235 170.355 ;
        RECT 46.525 170.185 46.695 170.355 ;
        RECT 46.985 170.185 47.155 170.355 ;
        RECT 47.445 170.185 47.615 170.355 ;
        RECT 47.905 170.185 48.075 170.355 ;
        RECT 48.365 170.185 48.535 170.355 ;
        RECT 48.825 170.185 48.995 170.355 ;
        RECT 49.285 170.185 49.455 170.355 ;
        RECT 49.745 170.185 49.915 170.355 ;
        RECT 50.205 170.185 50.375 170.355 ;
        RECT 50.665 170.185 50.835 170.355 ;
        RECT 51.125 170.185 51.295 170.355 ;
        RECT 51.585 170.185 51.755 170.355 ;
        RECT 52.045 170.185 52.215 170.355 ;
        RECT 52.505 170.185 52.675 170.355 ;
        RECT 52.965 170.185 53.135 170.355 ;
        RECT 53.425 170.185 53.595 170.355 ;
        RECT 53.885 170.185 54.055 170.355 ;
        RECT 54.345 170.185 54.515 170.355 ;
        RECT 54.805 170.185 54.975 170.355 ;
        RECT 55.265 170.185 55.435 170.355 ;
        RECT 55.725 170.185 55.895 170.355 ;
        RECT 56.185 170.185 56.355 170.355 ;
        RECT 56.645 170.185 56.815 170.355 ;
        RECT 57.105 170.185 57.275 170.355 ;
        RECT 57.565 170.185 57.735 170.355 ;
        RECT 58.025 170.185 58.195 170.355 ;
        RECT 58.485 170.185 58.655 170.355 ;
        RECT 58.945 170.185 59.115 170.355 ;
        RECT 59.405 170.185 59.575 170.355 ;
        RECT 59.865 170.185 60.035 170.355 ;
        RECT 60.325 170.185 60.495 170.355 ;
        RECT 60.785 170.185 60.955 170.355 ;
        RECT 61.245 170.185 61.415 170.355 ;
        RECT 61.705 170.185 61.875 170.355 ;
        RECT 62.165 170.185 62.335 170.355 ;
        RECT 62.625 170.185 62.795 170.355 ;
        RECT 63.085 170.185 63.255 170.355 ;
        RECT 63.545 170.185 63.715 170.355 ;
        RECT 64.005 170.185 64.175 170.355 ;
        RECT 64.465 170.185 64.635 170.355 ;
        RECT 64.925 170.185 65.095 170.355 ;
        RECT 65.385 170.185 65.555 170.355 ;
        RECT 65.845 170.185 66.015 170.355 ;
        RECT 66.305 170.185 66.475 170.355 ;
        RECT 66.765 170.185 66.935 170.355 ;
        RECT 67.225 170.185 67.395 170.355 ;
        RECT 67.685 170.185 67.855 170.355 ;
        RECT 68.145 170.185 68.315 170.355 ;
        RECT 68.605 170.185 68.775 170.355 ;
        RECT 69.065 170.185 69.235 170.355 ;
        RECT 69.525 170.185 69.695 170.355 ;
        RECT 69.985 170.185 70.155 170.355 ;
        RECT 70.445 170.185 70.615 170.355 ;
        RECT 70.905 170.185 71.075 170.355 ;
        RECT 71.365 170.185 71.535 170.355 ;
        RECT 71.825 170.185 71.995 170.355 ;
        RECT 72.285 170.185 72.455 170.355 ;
        RECT 72.745 170.185 72.915 170.355 ;
        RECT 73.205 170.185 73.375 170.355 ;
        RECT 73.665 170.185 73.835 170.355 ;
        RECT 74.125 170.185 74.295 170.355 ;
        RECT 74.585 170.185 74.755 170.355 ;
        RECT 75.045 170.185 75.215 170.355 ;
        RECT 75.505 170.185 75.675 170.355 ;
        RECT 75.965 170.185 76.135 170.355 ;
        RECT 76.425 170.185 76.595 170.355 ;
        RECT 76.885 170.185 77.055 170.355 ;
        RECT 77.345 170.185 77.515 170.355 ;
        RECT 77.805 170.185 77.975 170.355 ;
        RECT 78.265 170.185 78.435 170.355 ;
        RECT 78.725 170.185 78.895 170.355 ;
        RECT 79.185 170.185 79.355 170.355 ;
        RECT 79.645 170.185 79.815 170.355 ;
        RECT 80.105 170.185 80.275 170.355 ;
        RECT 80.565 170.185 80.735 170.355 ;
        RECT 81.025 170.185 81.195 170.355 ;
        RECT 81.485 170.185 81.655 170.355 ;
        RECT 81.945 170.185 82.115 170.355 ;
        RECT 82.405 170.185 82.575 170.355 ;
        RECT 82.865 170.185 83.035 170.355 ;
        RECT 83.325 170.185 83.495 170.355 ;
        RECT 83.785 170.185 83.955 170.355 ;
        RECT 84.245 170.185 84.415 170.355 ;
        RECT 84.705 170.185 84.875 170.355 ;
        RECT 85.165 170.185 85.335 170.355 ;
        RECT 85.625 170.185 85.795 170.355 ;
        RECT 86.085 170.185 86.255 170.355 ;
        RECT 86.545 170.185 86.715 170.355 ;
        RECT 87.005 170.185 87.175 170.355 ;
        RECT 87.465 170.185 87.635 170.355 ;
        RECT 87.925 170.185 88.095 170.355 ;
        RECT 88.385 170.185 88.555 170.355 ;
        RECT 88.845 170.185 89.015 170.355 ;
        RECT 89.305 170.185 89.475 170.355 ;
        RECT 89.765 170.185 89.935 170.355 ;
        RECT 90.225 170.185 90.395 170.355 ;
        RECT 90.685 170.185 90.855 170.355 ;
        RECT 91.145 170.185 91.315 170.355 ;
        RECT 91.605 170.185 91.775 170.355 ;
        RECT 92.065 170.185 92.235 170.355 ;
        RECT 92.525 170.185 92.695 170.355 ;
        RECT 92.985 170.185 93.155 170.355 ;
        RECT 93.445 170.185 93.615 170.355 ;
        RECT 93.905 170.185 94.075 170.355 ;
        RECT 94.365 170.185 94.535 170.355 ;
        RECT 94.825 170.185 94.995 170.355 ;
        RECT 95.285 170.185 95.455 170.355 ;
        RECT 95.745 170.185 95.915 170.355 ;
        RECT 96.205 170.185 96.375 170.355 ;
        RECT 96.665 170.185 96.835 170.355 ;
        RECT 97.125 170.185 97.295 170.355 ;
        RECT 97.585 170.185 97.755 170.355 ;
        RECT 98.045 170.185 98.215 170.355 ;
        RECT 98.505 170.185 98.675 170.355 ;
        RECT 98.965 170.185 99.135 170.355 ;
        RECT 99.425 170.185 99.595 170.355 ;
        RECT 99.885 170.185 100.055 170.355 ;
        RECT 100.345 170.185 100.515 170.355 ;
        RECT 100.805 170.185 100.975 170.355 ;
        RECT 101.265 170.185 101.435 170.355 ;
        RECT 101.725 170.185 101.895 170.355 ;
        RECT 102.185 170.185 102.355 170.355 ;
        RECT 102.645 170.185 102.815 170.355 ;
        RECT 103.105 170.185 103.275 170.355 ;
        RECT 103.565 170.185 103.735 170.355 ;
        RECT 104.025 170.185 104.195 170.355 ;
        RECT 104.485 170.185 104.655 170.355 ;
        RECT 104.945 170.185 105.115 170.355 ;
        RECT 105.405 170.185 105.575 170.355 ;
        RECT 105.865 170.185 106.035 170.355 ;
        RECT 106.325 170.185 106.495 170.355 ;
        RECT 106.785 170.185 106.955 170.355 ;
        RECT 107.245 170.185 107.415 170.355 ;
        RECT 107.705 170.185 107.875 170.355 ;
        RECT 108.165 170.185 108.335 170.355 ;
        RECT 108.625 170.185 108.795 170.355 ;
        RECT 109.085 170.185 109.255 170.355 ;
        RECT 109.545 170.185 109.715 170.355 ;
        RECT 110.005 170.185 110.175 170.355 ;
        RECT 110.465 170.185 110.635 170.355 ;
        RECT 110.925 170.185 111.095 170.355 ;
        RECT 111.385 170.185 111.555 170.355 ;
        RECT 111.845 170.185 112.015 170.355 ;
        RECT 112.305 170.185 112.475 170.355 ;
        RECT 112.765 170.185 112.935 170.355 ;
        RECT 113.225 170.185 113.395 170.355 ;
        RECT 113.685 170.185 113.855 170.355 ;
        RECT 114.145 170.185 114.315 170.355 ;
        RECT 114.605 170.185 114.775 170.355 ;
        RECT 115.065 170.185 115.235 170.355 ;
        RECT 115.525 170.185 115.695 170.355 ;
        RECT 41.925 164.745 42.095 164.915 ;
        RECT 42.385 164.745 42.555 164.915 ;
        RECT 42.845 164.745 43.015 164.915 ;
        RECT 43.305 164.745 43.475 164.915 ;
        RECT 43.765 164.745 43.935 164.915 ;
        RECT 44.225 164.745 44.395 164.915 ;
        RECT 44.685 164.745 44.855 164.915 ;
        RECT 45.145 164.745 45.315 164.915 ;
        RECT 45.605 164.745 45.775 164.915 ;
        RECT 46.065 164.745 46.235 164.915 ;
        RECT 46.525 164.745 46.695 164.915 ;
        RECT 46.985 164.745 47.155 164.915 ;
        RECT 47.445 164.745 47.615 164.915 ;
        RECT 47.905 164.745 48.075 164.915 ;
        RECT 48.365 164.745 48.535 164.915 ;
        RECT 48.825 164.745 48.995 164.915 ;
        RECT 49.285 164.745 49.455 164.915 ;
        RECT 49.745 164.745 49.915 164.915 ;
        RECT 50.205 164.745 50.375 164.915 ;
        RECT 50.665 164.745 50.835 164.915 ;
        RECT 51.125 164.745 51.295 164.915 ;
        RECT 51.585 164.745 51.755 164.915 ;
        RECT 52.045 164.745 52.215 164.915 ;
        RECT 52.505 164.745 52.675 164.915 ;
        RECT 52.965 164.745 53.135 164.915 ;
        RECT 53.425 164.745 53.595 164.915 ;
        RECT 53.885 164.745 54.055 164.915 ;
        RECT 54.345 164.745 54.515 164.915 ;
        RECT 54.805 164.745 54.975 164.915 ;
        RECT 55.265 164.745 55.435 164.915 ;
        RECT 55.725 164.745 55.895 164.915 ;
        RECT 56.185 164.745 56.355 164.915 ;
        RECT 56.645 164.745 56.815 164.915 ;
        RECT 57.105 164.745 57.275 164.915 ;
        RECT 57.565 164.745 57.735 164.915 ;
        RECT 58.025 164.745 58.195 164.915 ;
        RECT 58.485 164.745 58.655 164.915 ;
        RECT 58.945 164.745 59.115 164.915 ;
        RECT 59.405 164.745 59.575 164.915 ;
        RECT 59.865 164.745 60.035 164.915 ;
        RECT 60.325 164.745 60.495 164.915 ;
        RECT 60.785 164.745 60.955 164.915 ;
        RECT 61.245 164.745 61.415 164.915 ;
        RECT 61.705 164.745 61.875 164.915 ;
        RECT 62.165 164.745 62.335 164.915 ;
        RECT 62.625 164.745 62.795 164.915 ;
        RECT 63.085 164.745 63.255 164.915 ;
        RECT 63.545 164.745 63.715 164.915 ;
        RECT 64.005 164.745 64.175 164.915 ;
        RECT 64.465 164.745 64.635 164.915 ;
        RECT 64.925 164.745 65.095 164.915 ;
        RECT 65.385 164.745 65.555 164.915 ;
        RECT 65.845 164.745 66.015 164.915 ;
        RECT 66.305 164.745 66.475 164.915 ;
        RECT 66.765 164.745 66.935 164.915 ;
        RECT 67.225 164.745 67.395 164.915 ;
        RECT 67.685 164.745 67.855 164.915 ;
        RECT 68.145 164.745 68.315 164.915 ;
        RECT 68.605 164.745 68.775 164.915 ;
        RECT 69.065 164.745 69.235 164.915 ;
        RECT 69.525 164.745 69.695 164.915 ;
        RECT 69.985 164.745 70.155 164.915 ;
        RECT 70.445 164.745 70.615 164.915 ;
        RECT 70.905 164.745 71.075 164.915 ;
        RECT 71.365 164.745 71.535 164.915 ;
        RECT 71.825 164.745 71.995 164.915 ;
        RECT 72.285 164.745 72.455 164.915 ;
        RECT 72.745 164.745 72.915 164.915 ;
        RECT 73.205 164.745 73.375 164.915 ;
        RECT 73.665 164.745 73.835 164.915 ;
        RECT 74.125 164.745 74.295 164.915 ;
        RECT 74.585 164.745 74.755 164.915 ;
        RECT 75.045 164.745 75.215 164.915 ;
        RECT 75.505 164.745 75.675 164.915 ;
        RECT 75.965 164.745 76.135 164.915 ;
        RECT 76.425 164.745 76.595 164.915 ;
        RECT 76.885 164.745 77.055 164.915 ;
        RECT 77.345 164.745 77.515 164.915 ;
        RECT 77.805 164.745 77.975 164.915 ;
        RECT 78.265 164.745 78.435 164.915 ;
        RECT 78.725 164.745 78.895 164.915 ;
        RECT 79.185 164.745 79.355 164.915 ;
        RECT 79.645 164.745 79.815 164.915 ;
        RECT 80.105 164.745 80.275 164.915 ;
        RECT 80.565 164.745 80.735 164.915 ;
        RECT 81.025 164.745 81.195 164.915 ;
        RECT 81.485 164.745 81.655 164.915 ;
        RECT 81.945 164.745 82.115 164.915 ;
        RECT 82.405 164.745 82.575 164.915 ;
        RECT 82.865 164.745 83.035 164.915 ;
        RECT 83.325 164.745 83.495 164.915 ;
        RECT 83.785 164.745 83.955 164.915 ;
        RECT 84.245 164.745 84.415 164.915 ;
        RECT 84.705 164.745 84.875 164.915 ;
        RECT 85.165 164.745 85.335 164.915 ;
        RECT 85.625 164.745 85.795 164.915 ;
        RECT 86.085 164.745 86.255 164.915 ;
        RECT 86.545 164.745 86.715 164.915 ;
        RECT 87.005 164.745 87.175 164.915 ;
        RECT 87.465 164.745 87.635 164.915 ;
        RECT 87.925 164.745 88.095 164.915 ;
        RECT 88.385 164.745 88.555 164.915 ;
        RECT 88.845 164.745 89.015 164.915 ;
        RECT 89.305 164.745 89.475 164.915 ;
        RECT 89.765 164.745 89.935 164.915 ;
        RECT 90.225 164.745 90.395 164.915 ;
        RECT 90.685 164.745 90.855 164.915 ;
        RECT 91.145 164.745 91.315 164.915 ;
        RECT 91.605 164.745 91.775 164.915 ;
        RECT 92.065 164.745 92.235 164.915 ;
        RECT 92.525 164.745 92.695 164.915 ;
        RECT 92.985 164.745 93.155 164.915 ;
        RECT 93.445 164.745 93.615 164.915 ;
        RECT 93.905 164.745 94.075 164.915 ;
        RECT 94.365 164.745 94.535 164.915 ;
        RECT 94.825 164.745 94.995 164.915 ;
        RECT 95.285 164.745 95.455 164.915 ;
        RECT 95.745 164.745 95.915 164.915 ;
        RECT 96.205 164.745 96.375 164.915 ;
        RECT 96.665 164.745 96.835 164.915 ;
        RECT 97.125 164.745 97.295 164.915 ;
        RECT 97.585 164.745 97.755 164.915 ;
        RECT 98.045 164.745 98.215 164.915 ;
        RECT 98.505 164.745 98.675 164.915 ;
        RECT 98.965 164.745 99.135 164.915 ;
        RECT 99.425 164.745 99.595 164.915 ;
        RECT 99.885 164.745 100.055 164.915 ;
        RECT 100.345 164.745 100.515 164.915 ;
        RECT 100.805 164.745 100.975 164.915 ;
        RECT 101.265 164.745 101.435 164.915 ;
        RECT 101.725 164.745 101.895 164.915 ;
        RECT 102.185 164.745 102.355 164.915 ;
        RECT 102.645 164.745 102.815 164.915 ;
        RECT 103.105 164.745 103.275 164.915 ;
        RECT 103.565 164.745 103.735 164.915 ;
        RECT 104.025 164.745 104.195 164.915 ;
        RECT 104.485 164.745 104.655 164.915 ;
        RECT 104.945 164.745 105.115 164.915 ;
        RECT 105.405 164.745 105.575 164.915 ;
        RECT 105.865 164.745 106.035 164.915 ;
        RECT 106.325 164.745 106.495 164.915 ;
        RECT 106.785 164.745 106.955 164.915 ;
        RECT 107.245 164.745 107.415 164.915 ;
        RECT 107.705 164.745 107.875 164.915 ;
        RECT 108.165 164.745 108.335 164.915 ;
        RECT 108.625 164.745 108.795 164.915 ;
        RECT 109.085 164.745 109.255 164.915 ;
        RECT 109.545 164.745 109.715 164.915 ;
        RECT 110.005 164.745 110.175 164.915 ;
        RECT 110.465 164.745 110.635 164.915 ;
        RECT 110.925 164.745 111.095 164.915 ;
        RECT 111.385 164.745 111.555 164.915 ;
        RECT 111.845 164.745 112.015 164.915 ;
        RECT 112.305 164.745 112.475 164.915 ;
        RECT 112.765 164.745 112.935 164.915 ;
        RECT 113.225 164.745 113.395 164.915 ;
        RECT 113.685 164.745 113.855 164.915 ;
        RECT 114.145 164.745 114.315 164.915 ;
        RECT 114.605 164.745 114.775 164.915 ;
        RECT 115.065 164.745 115.235 164.915 ;
        RECT 115.525 164.745 115.695 164.915 ;
        RECT 41.925 159.305 42.095 159.475 ;
        RECT 42.385 159.305 42.555 159.475 ;
        RECT 42.845 159.305 43.015 159.475 ;
        RECT 43.305 159.305 43.475 159.475 ;
        RECT 43.765 159.305 43.935 159.475 ;
        RECT 44.225 159.305 44.395 159.475 ;
        RECT 44.685 159.305 44.855 159.475 ;
        RECT 45.145 159.305 45.315 159.475 ;
        RECT 45.605 159.305 45.775 159.475 ;
        RECT 46.065 159.305 46.235 159.475 ;
        RECT 46.525 159.305 46.695 159.475 ;
        RECT 46.985 159.305 47.155 159.475 ;
        RECT 47.445 159.305 47.615 159.475 ;
        RECT 47.905 159.305 48.075 159.475 ;
        RECT 48.365 159.305 48.535 159.475 ;
        RECT 48.825 159.305 48.995 159.475 ;
        RECT 49.285 159.305 49.455 159.475 ;
        RECT 49.745 159.305 49.915 159.475 ;
        RECT 50.205 159.305 50.375 159.475 ;
        RECT 50.665 159.305 50.835 159.475 ;
        RECT 51.125 159.305 51.295 159.475 ;
        RECT 51.585 159.305 51.755 159.475 ;
        RECT 52.045 159.305 52.215 159.475 ;
        RECT 52.505 159.305 52.675 159.475 ;
        RECT 52.965 159.305 53.135 159.475 ;
        RECT 53.425 159.305 53.595 159.475 ;
        RECT 53.885 159.305 54.055 159.475 ;
        RECT 54.345 159.305 54.515 159.475 ;
        RECT 54.805 159.305 54.975 159.475 ;
        RECT 55.265 159.305 55.435 159.475 ;
        RECT 55.725 159.305 55.895 159.475 ;
        RECT 56.185 159.305 56.355 159.475 ;
        RECT 56.645 159.305 56.815 159.475 ;
        RECT 57.105 159.305 57.275 159.475 ;
        RECT 57.565 159.305 57.735 159.475 ;
        RECT 58.025 159.305 58.195 159.475 ;
        RECT 58.485 159.305 58.655 159.475 ;
        RECT 58.945 159.305 59.115 159.475 ;
        RECT 59.405 159.305 59.575 159.475 ;
        RECT 59.865 159.305 60.035 159.475 ;
        RECT 60.325 159.305 60.495 159.475 ;
        RECT 60.785 159.305 60.955 159.475 ;
        RECT 61.245 159.305 61.415 159.475 ;
        RECT 61.705 159.305 61.875 159.475 ;
        RECT 62.165 159.305 62.335 159.475 ;
        RECT 62.625 159.305 62.795 159.475 ;
        RECT 63.085 159.305 63.255 159.475 ;
        RECT 63.545 159.305 63.715 159.475 ;
        RECT 64.005 159.305 64.175 159.475 ;
        RECT 64.465 159.305 64.635 159.475 ;
        RECT 64.925 159.305 65.095 159.475 ;
        RECT 65.385 159.305 65.555 159.475 ;
        RECT 65.845 159.305 66.015 159.475 ;
        RECT 66.305 159.305 66.475 159.475 ;
        RECT 66.765 159.305 66.935 159.475 ;
        RECT 67.225 159.305 67.395 159.475 ;
        RECT 67.685 159.305 67.855 159.475 ;
        RECT 68.145 159.305 68.315 159.475 ;
        RECT 68.605 159.305 68.775 159.475 ;
        RECT 69.065 159.305 69.235 159.475 ;
        RECT 69.525 159.305 69.695 159.475 ;
        RECT 69.985 159.305 70.155 159.475 ;
        RECT 70.445 159.305 70.615 159.475 ;
        RECT 70.905 159.305 71.075 159.475 ;
        RECT 71.365 159.305 71.535 159.475 ;
        RECT 71.825 159.305 71.995 159.475 ;
        RECT 72.285 159.305 72.455 159.475 ;
        RECT 72.745 159.305 72.915 159.475 ;
        RECT 73.205 159.305 73.375 159.475 ;
        RECT 73.665 159.305 73.835 159.475 ;
        RECT 74.125 159.305 74.295 159.475 ;
        RECT 74.585 159.305 74.755 159.475 ;
        RECT 75.045 159.305 75.215 159.475 ;
        RECT 75.505 159.305 75.675 159.475 ;
        RECT 75.965 159.305 76.135 159.475 ;
        RECT 76.425 159.305 76.595 159.475 ;
        RECT 76.885 159.305 77.055 159.475 ;
        RECT 77.345 159.305 77.515 159.475 ;
        RECT 77.805 159.305 77.975 159.475 ;
        RECT 78.265 159.305 78.435 159.475 ;
        RECT 78.725 159.305 78.895 159.475 ;
        RECT 79.185 159.305 79.355 159.475 ;
        RECT 79.645 159.305 79.815 159.475 ;
        RECT 80.105 159.305 80.275 159.475 ;
        RECT 80.565 159.305 80.735 159.475 ;
        RECT 81.025 159.305 81.195 159.475 ;
        RECT 81.485 159.305 81.655 159.475 ;
        RECT 81.945 159.305 82.115 159.475 ;
        RECT 82.405 159.305 82.575 159.475 ;
        RECT 82.865 159.305 83.035 159.475 ;
        RECT 83.325 159.305 83.495 159.475 ;
        RECT 83.785 159.305 83.955 159.475 ;
        RECT 84.245 159.305 84.415 159.475 ;
        RECT 84.705 159.305 84.875 159.475 ;
        RECT 85.165 159.305 85.335 159.475 ;
        RECT 85.625 159.305 85.795 159.475 ;
        RECT 86.085 159.305 86.255 159.475 ;
        RECT 86.545 159.305 86.715 159.475 ;
        RECT 87.005 159.305 87.175 159.475 ;
        RECT 87.465 159.305 87.635 159.475 ;
        RECT 87.925 159.305 88.095 159.475 ;
        RECT 88.385 159.305 88.555 159.475 ;
        RECT 88.845 159.305 89.015 159.475 ;
        RECT 89.305 159.305 89.475 159.475 ;
        RECT 89.765 159.305 89.935 159.475 ;
        RECT 90.225 159.305 90.395 159.475 ;
        RECT 90.685 159.305 90.855 159.475 ;
        RECT 91.145 159.305 91.315 159.475 ;
        RECT 91.605 159.305 91.775 159.475 ;
        RECT 92.065 159.305 92.235 159.475 ;
        RECT 92.525 159.305 92.695 159.475 ;
        RECT 92.985 159.305 93.155 159.475 ;
        RECT 93.445 159.305 93.615 159.475 ;
        RECT 93.905 159.305 94.075 159.475 ;
        RECT 94.365 159.305 94.535 159.475 ;
        RECT 94.825 159.305 94.995 159.475 ;
        RECT 95.285 159.305 95.455 159.475 ;
        RECT 95.745 159.305 95.915 159.475 ;
        RECT 96.205 159.305 96.375 159.475 ;
        RECT 96.665 159.305 96.835 159.475 ;
        RECT 97.125 159.305 97.295 159.475 ;
        RECT 97.585 159.305 97.755 159.475 ;
        RECT 98.045 159.305 98.215 159.475 ;
        RECT 98.505 159.305 98.675 159.475 ;
        RECT 98.965 159.305 99.135 159.475 ;
        RECT 99.425 159.305 99.595 159.475 ;
        RECT 99.885 159.305 100.055 159.475 ;
        RECT 100.345 159.305 100.515 159.475 ;
        RECT 100.805 159.305 100.975 159.475 ;
        RECT 101.265 159.305 101.435 159.475 ;
        RECT 101.725 159.305 101.895 159.475 ;
        RECT 102.185 159.305 102.355 159.475 ;
        RECT 102.645 159.305 102.815 159.475 ;
        RECT 103.105 159.305 103.275 159.475 ;
        RECT 103.565 159.305 103.735 159.475 ;
        RECT 104.025 159.305 104.195 159.475 ;
        RECT 104.485 159.305 104.655 159.475 ;
        RECT 104.945 159.305 105.115 159.475 ;
        RECT 105.405 159.305 105.575 159.475 ;
        RECT 105.865 159.305 106.035 159.475 ;
        RECT 106.325 159.305 106.495 159.475 ;
        RECT 106.785 159.305 106.955 159.475 ;
        RECT 107.245 159.305 107.415 159.475 ;
        RECT 107.705 159.305 107.875 159.475 ;
        RECT 108.165 159.305 108.335 159.475 ;
        RECT 108.625 159.305 108.795 159.475 ;
        RECT 109.085 159.305 109.255 159.475 ;
        RECT 109.545 159.305 109.715 159.475 ;
        RECT 110.005 159.305 110.175 159.475 ;
        RECT 110.465 159.305 110.635 159.475 ;
        RECT 110.925 159.305 111.095 159.475 ;
        RECT 111.385 159.305 111.555 159.475 ;
        RECT 111.845 159.305 112.015 159.475 ;
        RECT 112.305 159.305 112.475 159.475 ;
        RECT 112.765 159.305 112.935 159.475 ;
        RECT 113.225 159.305 113.395 159.475 ;
        RECT 113.685 159.305 113.855 159.475 ;
        RECT 114.145 159.305 114.315 159.475 ;
        RECT 114.605 159.305 114.775 159.475 ;
        RECT 115.065 159.305 115.235 159.475 ;
        RECT 115.525 159.305 115.695 159.475 ;
        RECT 59.470 119.540 59.640 120.420 ;
        RECT 60.870 119.540 61.040 120.420 ;
        RECT 58.145 119.085 58.315 119.255 ;
        RECT 67.700 117.350 67.870 121.230 ;
        RECT 68.290 117.350 68.460 121.230 ;
        RECT 70.170 117.350 70.340 121.230 ;
        RECT 72.050 117.350 72.220 121.230 ;
        RECT 76.620 119.445 76.810 121.430 ;
        RECT 82.130 119.540 82.300 120.420 ;
        RECT 83.530 119.540 83.700 120.420 ;
        RECT 80.805 119.085 80.975 119.255 ;
        RECT 90.360 117.350 90.530 121.230 ;
        RECT 90.950 117.350 91.120 121.230 ;
        RECT 92.830 117.350 93.000 121.230 ;
        RECT 94.710 117.350 94.880 121.230 ;
        RECT 99.280 119.445 99.470 121.430 ;
        RECT 104.790 119.540 104.960 120.420 ;
        RECT 106.190 119.540 106.360 120.420 ;
        RECT 103.465 119.085 103.635 119.255 ;
        RECT 113.020 117.350 113.190 121.230 ;
        RECT 113.610 117.350 113.780 121.230 ;
        RECT 115.490 117.350 115.660 121.230 ;
        RECT 117.370 117.350 117.540 121.230 ;
        RECT 121.940 119.445 122.130 121.430 ;
        RECT 67.700 112.170 67.870 116.050 ;
        RECT 68.290 112.170 68.460 116.050 ;
        RECT 70.170 112.170 70.340 116.050 ;
        RECT 72.050 112.170 72.220 116.050 ;
        RECT 90.360 112.170 90.530 116.050 ;
        RECT 90.950 112.170 91.120 116.050 ;
        RECT 92.830 112.170 93.000 116.050 ;
        RECT 94.710 112.170 94.880 116.050 ;
        RECT 113.020 112.170 113.190 116.050 ;
        RECT 113.610 112.170 113.780 116.050 ;
        RECT 115.490 112.170 115.660 116.050 ;
        RECT 117.370 112.170 117.540 116.050 ;
        RECT 64.190 111.480 64.400 111.690 ;
        RECT 66.070 111.480 66.280 111.690 ;
        RECT 67.950 111.480 68.160 111.690 ;
        RECT 69.830 111.480 70.040 111.690 ;
        RECT 71.710 111.480 71.920 111.690 ;
        RECT 86.850 111.480 87.060 111.690 ;
        RECT 88.730 111.480 88.940 111.690 ;
        RECT 90.610 111.480 90.820 111.690 ;
        RECT 92.490 111.480 92.700 111.690 ;
        RECT 94.370 111.480 94.580 111.690 ;
        RECT 109.510 111.480 109.720 111.690 ;
        RECT 111.390 111.480 111.600 111.690 ;
        RECT 113.270 111.480 113.480 111.690 ;
        RECT 115.150 111.480 115.360 111.690 ;
        RECT 117.030 111.480 117.240 111.690 ;
        RECT 56.300 107.365 56.490 109.350 ;
        RECT 36.810 102.200 36.980 103.080 ;
        RECT 38.210 102.200 38.380 103.080 ;
        RECT 35.485 101.745 35.655 101.915 ;
        RECT 45.040 100.010 45.210 103.890 ;
        RECT 45.630 100.010 45.800 103.890 ;
        RECT 47.510 100.010 47.680 103.890 ;
        RECT 49.390 100.010 49.560 103.890 ;
        RECT 53.960 102.105 54.150 104.090 ;
        RECT 59.470 102.200 59.640 103.080 ;
        RECT 60.870 102.200 61.040 103.080 ;
        RECT 58.145 101.745 58.315 101.915 ;
        RECT 67.700 100.010 67.870 103.890 ;
        RECT 68.290 100.010 68.460 103.890 ;
        RECT 70.170 100.010 70.340 103.890 ;
        RECT 72.050 100.010 72.220 103.890 ;
        RECT 76.620 102.105 76.810 104.090 ;
        RECT 82.130 102.200 82.300 103.080 ;
        RECT 83.530 102.200 83.700 103.080 ;
        RECT 80.805 101.745 80.975 101.915 ;
        RECT 90.360 100.010 90.530 103.890 ;
        RECT 90.950 100.010 91.120 103.890 ;
        RECT 92.830 100.010 93.000 103.890 ;
        RECT 94.710 100.010 94.880 103.890 ;
        RECT 99.280 102.105 99.470 104.090 ;
        RECT 104.790 102.200 104.960 103.080 ;
        RECT 106.190 102.200 106.360 103.080 ;
        RECT 103.465 101.745 103.635 101.915 ;
        RECT 113.020 100.010 113.190 103.890 ;
        RECT 113.610 100.010 113.780 103.890 ;
        RECT 115.490 100.010 115.660 103.890 ;
        RECT 117.370 100.010 117.540 103.890 ;
        RECT 121.940 102.105 122.130 104.090 ;
        RECT 45.040 94.830 45.210 98.710 ;
        RECT 45.630 94.830 45.800 98.710 ;
        RECT 47.510 94.830 47.680 98.710 ;
        RECT 49.390 94.830 49.560 98.710 ;
        RECT 67.700 94.830 67.870 98.710 ;
        RECT 68.290 94.830 68.460 98.710 ;
        RECT 70.170 94.830 70.340 98.710 ;
        RECT 72.050 94.830 72.220 98.710 ;
        RECT 90.360 94.830 90.530 98.710 ;
        RECT 90.950 94.830 91.120 98.710 ;
        RECT 92.830 94.830 93.000 98.710 ;
        RECT 94.710 94.830 94.880 98.710 ;
        RECT 113.020 94.830 113.190 98.710 ;
        RECT 113.610 94.830 113.780 98.710 ;
        RECT 115.490 94.830 115.660 98.710 ;
        RECT 117.370 94.830 117.540 98.710 ;
        RECT 41.530 94.140 41.740 94.350 ;
        RECT 43.410 94.140 43.620 94.350 ;
        RECT 45.290 94.140 45.500 94.350 ;
        RECT 47.170 94.140 47.380 94.350 ;
        RECT 49.050 94.140 49.260 94.350 ;
        RECT 64.190 94.140 64.400 94.350 ;
        RECT 66.070 94.140 66.280 94.350 ;
        RECT 67.950 94.140 68.160 94.350 ;
        RECT 69.830 94.140 70.040 94.350 ;
        RECT 71.710 94.140 71.920 94.350 ;
        RECT 86.850 94.140 87.060 94.350 ;
        RECT 88.730 94.140 88.940 94.350 ;
        RECT 90.610 94.140 90.820 94.350 ;
        RECT 92.490 94.140 92.700 94.350 ;
        RECT 94.370 94.140 94.580 94.350 ;
        RECT 109.510 94.140 109.720 94.350 ;
        RECT 111.390 94.140 111.600 94.350 ;
        RECT 113.270 94.140 113.480 94.350 ;
        RECT 115.150 94.140 115.360 94.350 ;
        RECT 117.030 94.140 117.240 94.350 ;
        RECT 36.810 84.860 36.980 85.740 ;
        RECT 38.210 84.860 38.380 85.740 ;
        RECT 35.485 84.405 35.655 84.575 ;
        RECT 45.040 82.670 45.210 86.550 ;
        RECT 45.630 82.670 45.800 86.550 ;
        RECT 47.510 82.670 47.680 86.550 ;
        RECT 49.390 82.670 49.560 86.550 ;
        RECT 53.960 84.765 54.150 86.750 ;
        RECT 59.470 84.860 59.640 85.740 ;
        RECT 60.870 84.860 61.040 85.740 ;
        RECT 58.145 84.405 58.315 84.575 ;
        RECT 67.700 82.670 67.870 86.550 ;
        RECT 68.290 82.670 68.460 86.550 ;
        RECT 70.170 82.670 70.340 86.550 ;
        RECT 72.050 82.670 72.220 86.550 ;
        RECT 76.620 84.765 76.810 86.750 ;
        RECT 82.130 84.860 82.300 85.740 ;
        RECT 83.530 84.860 83.700 85.740 ;
        RECT 80.805 84.405 80.975 84.575 ;
        RECT 90.360 82.670 90.530 86.550 ;
        RECT 90.950 82.670 91.120 86.550 ;
        RECT 92.830 82.670 93.000 86.550 ;
        RECT 94.710 82.670 94.880 86.550 ;
        RECT 99.280 84.765 99.470 86.750 ;
        RECT 104.790 84.860 104.960 85.740 ;
        RECT 106.190 84.860 106.360 85.740 ;
        RECT 103.465 84.405 103.635 84.575 ;
        RECT 113.020 82.670 113.190 86.550 ;
        RECT 113.610 82.670 113.780 86.550 ;
        RECT 115.490 82.670 115.660 86.550 ;
        RECT 117.370 82.670 117.540 86.550 ;
        RECT 121.940 84.765 122.130 86.750 ;
        RECT 45.040 77.490 45.210 81.370 ;
        RECT 45.630 77.490 45.800 81.370 ;
        RECT 47.510 77.490 47.680 81.370 ;
        RECT 49.390 77.490 49.560 81.370 ;
        RECT 67.700 77.490 67.870 81.370 ;
        RECT 68.290 77.490 68.460 81.370 ;
        RECT 70.170 77.490 70.340 81.370 ;
        RECT 72.050 77.490 72.220 81.370 ;
        RECT 90.360 77.490 90.530 81.370 ;
        RECT 90.950 77.490 91.120 81.370 ;
        RECT 92.830 77.490 93.000 81.370 ;
        RECT 94.710 77.490 94.880 81.370 ;
        RECT 113.020 77.490 113.190 81.370 ;
        RECT 113.610 77.490 113.780 81.370 ;
        RECT 115.490 77.490 115.660 81.370 ;
        RECT 117.370 77.490 117.540 81.370 ;
        RECT 41.530 76.800 41.740 77.010 ;
        RECT 43.410 76.800 43.620 77.010 ;
        RECT 45.290 76.800 45.500 77.010 ;
        RECT 47.170 76.800 47.380 77.010 ;
        RECT 49.050 76.800 49.260 77.010 ;
        RECT 64.190 76.800 64.400 77.010 ;
        RECT 66.070 76.800 66.280 77.010 ;
        RECT 67.950 76.800 68.160 77.010 ;
        RECT 69.830 76.800 70.040 77.010 ;
        RECT 71.710 76.800 71.920 77.010 ;
        RECT 86.850 76.800 87.060 77.010 ;
        RECT 88.730 76.800 88.940 77.010 ;
        RECT 90.610 76.800 90.820 77.010 ;
        RECT 92.490 76.800 92.700 77.010 ;
        RECT 94.370 76.800 94.580 77.010 ;
        RECT 109.510 76.800 109.720 77.010 ;
        RECT 111.390 76.800 111.600 77.010 ;
        RECT 113.270 76.800 113.480 77.010 ;
        RECT 115.150 76.800 115.360 77.010 ;
        RECT 117.030 76.800 117.240 77.010 ;
        RECT 36.810 67.520 36.980 68.400 ;
        RECT 38.210 67.520 38.380 68.400 ;
        RECT 35.485 67.065 35.655 67.235 ;
        RECT 45.040 65.330 45.210 69.210 ;
        RECT 45.630 65.330 45.800 69.210 ;
        RECT 47.510 65.330 47.680 69.210 ;
        RECT 49.390 65.330 49.560 69.210 ;
        RECT 53.960 67.425 54.150 69.410 ;
        RECT 59.470 67.520 59.640 68.400 ;
        RECT 60.870 67.520 61.040 68.400 ;
        RECT 58.145 67.065 58.315 67.235 ;
        RECT 67.700 65.330 67.870 69.210 ;
        RECT 68.290 65.330 68.460 69.210 ;
        RECT 70.170 65.330 70.340 69.210 ;
        RECT 72.050 65.330 72.220 69.210 ;
        RECT 76.620 67.425 76.810 69.410 ;
        RECT 82.130 67.520 82.300 68.400 ;
        RECT 83.530 67.520 83.700 68.400 ;
        RECT 80.805 67.065 80.975 67.235 ;
        RECT 90.360 65.330 90.530 69.210 ;
        RECT 90.950 65.330 91.120 69.210 ;
        RECT 92.830 65.330 93.000 69.210 ;
        RECT 94.710 65.330 94.880 69.210 ;
        RECT 99.280 67.425 99.470 69.410 ;
        RECT 104.790 67.520 104.960 68.400 ;
        RECT 106.190 67.520 106.360 68.400 ;
        RECT 103.465 67.065 103.635 67.235 ;
        RECT 113.020 65.330 113.190 69.210 ;
        RECT 113.610 65.330 113.780 69.210 ;
        RECT 115.490 65.330 115.660 69.210 ;
        RECT 117.370 65.330 117.540 69.210 ;
        RECT 121.940 67.425 122.130 69.410 ;
        RECT 45.040 60.150 45.210 64.030 ;
        RECT 45.630 60.150 45.800 64.030 ;
        RECT 47.510 60.150 47.680 64.030 ;
        RECT 49.390 60.150 49.560 64.030 ;
        RECT 67.700 60.150 67.870 64.030 ;
        RECT 68.290 60.150 68.460 64.030 ;
        RECT 70.170 60.150 70.340 64.030 ;
        RECT 72.050 60.150 72.220 64.030 ;
        RECT 90.360 60.150 90.530 64.030 ;
        RECT 90.950 60.150 91.120 64.030 ;
        RECT 92.830 60.150 93.000 64.030 ;
        RECT 94.710 60.150 94.880 64.030 ;
        RECT 113.020 60.150 113.190 64.030 ;
        RECT 113.610 60.150 113.780 64.030 ;
        RECT 115.490 60.150 115.660 64.030 ;
        RECT 117.370 60.150 117.540 64.030 ;
        RECT 41.530 59.460 41.740 59.670 ;
        RECT 43.410 59.460 43.620 59.670 ;
        RECT 45.290 59.460 45.500 59.670 ;
        RECT 47.170 59.460 47.380 59.670 ;
        RECT 49.050 59.460 49.260 59.670 ;
        RECT 64.190 59.460 64.400 59.670 ;
        RECT 66.070 59.460 66.280 59.670 ;
        RECT 67.950 59.460 68.160 59.670 ;
        RECT 69.830 59.460 70.040 59.670 ;
        RECT 71.710 59.460 71.920 59.670 ;
        RECT 86.850 59.460 87.060 59.670 ;
        RECT 88.730 59.460 88.940 59.670 ;
        RECT 90.610 59.460 90.820 59.670 ;
        RECT 92.490 59.460 92.700 59.670 ;
        RECT 94.370 59.460 94.580 59.670 ;
        RECT 109.510 59.460 109.720 59.670 ;
        RECT 111.390 59.460 111.600 59.670 ;
        RECT 113.270 59.460 113.480 59.670 ;
        RECT 115.150 59.460 115.360 59.670 ;
        RECT 117.030 59.460 117.240 59.670 ;
        RECT 45.040 47.330 45.210 51.210 ;
        RECT 45.630 47.330 45.800 51.210 ;
        RECT 47.510 47.330 47.680 51.210 ;
        RECT 49.390 47.330 49.560 51.210 ;
        RECT 53.960 49.425 54.150 51.410 ;
        RECT 67.700 47.330 67.870 51.210 ;
        RECT 68.290 47.330 68.460 51.210 ;
        RECT 70.170 47.330 70.340 51.210 ;
        RECT 72.050 47.330 72.220 51.210 ;
        RECT 76.620 49.425 76.810 51.410 ;
        RECT 90.360 47.330 90.530 51.210 ;
        RECT 90.950 47.330 91.120 51.210 ;
        RECT 92.830 47.330 93.000 51.210 ;
        RECT 94.710 47.330 94.880 51.210 ;
        RECT 99.280 49.425 99.470 51.410 ;
        RECT 113.020 47.330 113.190 51.210 ;
        RECT 113.610 47.330 113.780 51.210 ;
        RECT 115.490 47.330 115.660 51.210 ;
        RECT 117.370 47.330 117.540 51.210 ;
        RECT 121.940 49.425 122.130 51.410 ;
        RECT 45.040 42.150 45.210 46.030 ;
        RECT 45.630 42.150 45.800 46.030 ;
        RECT 47.510 42.150 47.680 46.030 ;
        RECT 49.390 42.150 49.560 46.030 ;
        RECT 67.700 42.150 67.870 46.030 ;
        RECT 68.290 42.150 68.460 46.030 ;
        RECT 70.170 42.150 70.340 46.030 ;
        RECT 72.050 42.150 72.220 46.030 ;
        RECT 90.360 42.150 90.530 46.030 ;
        RECT 90.950 42.150 91.120 46.030 ;
        RECT 92.830 42.150 93.000 46.030 ;
        RECT 94.710 42.150 94.880 46.030 ;
        RECT 113.020 42.150 113.190 46.030 ;
        RECT 113.610 42.150 113.780 46.030 ;
        RECT 115.490 42.150 115.660 46.030 ;
        RECT 117.370 42.150 117.540 46.030 ;
        RECT 41.530 41.460 41.740 41.670 ;
        RECT 43.410 41.460 43.620 41.670 ;
        RECT 45.290 41.460 45.500 41.670 ;
        RECT 47.170 41.460 47.380 41.670 ;
        RECT 49.050 41.460 49.260 41.670 ;
        RECT 64.190 41.460 64.400 41.670 ;
        RECT 66.070 41.460 66.280 41.670 ;
        RECT 67.950 41.460 68.160 41.670 ;
        RECT 69.830 41.460 70.040 41.670 ;
        RECT 71.710 41.460 71.920 41.670 ;
        RECT 86.850 41.460 87.060 41.670 ;
        RECT 88.730 41.460 88.940 41.670 ;
        RECT 90.610 41.460 90.820 41.670 ;
        RECT 92.490 41.460 92.700 41.670 ;
        RECT 94.370 41.460 94.580 41.670 ;
        RECT 109.510 41.460 109.720 41.670 ;
        RECT 111.390 41.460 111.600 41.670 ;
        RECT 113.270 41.460 113.480 41.670 ;
        RECT 115.150 41.460 115.360 41.670 ;
        RECT 117.030 41.460 117.240 41.670 ;
      LAYER met1 ;
        RECT 41.780 186.350 115.840 186.830 ;
        RECT 41.780 180.910 115.840 181.390 ;
        RECT 41.780 175.470 115.840 175.950 ;
        RECT 41.780 170.030 115.840 170.510 ;
        RECT 41.780 164.590 115.840 165.070 ;
        RECT 41.780 159.150 115.840 159.630 ;
        RECT 67.670 121.240 67.900 121.290 ;
        RECT 68.260 121.240 68.490 121.290 ;
        RECT 67.670 121.050 68.490 121.240 ;
        RECT 59.440 119.605 59.670 120.480 ;
        RECT 60.840 119.965 61.070 120.480 ;
        RECT 61.250 119.965 62.250 119.980 ;
        RECT 60.840 119.775 62.250 119.965 ;
        RECT 59.440 119.480 59.865 119.605 ;
        RECT 60.840 119.480 61.070 119.775 ;
        RECT 59.460 119.415 59.865 119.480 ;
        RECT 58.085 119.265 58.375 119.285 ;
        RECT 58.085 119.055 58.645 119.265 ;
        RECT 58.455 118.905 58.645 119.055 ;
        RECT 59.675 118.905 59.865 119.415 ;
        RECT 61.250 118.980 62.250 119.775 ;
        RECT 61.250 118.905 61.440 118.980 ;
        RECT 58.455 118.715 61.440 118.905 ;
        RECT 67.670 117.540 67.900 121.050 ;
        RECT 68.260 117.540 68.490 121.050 ;
        RECT 67.670 117.290 68.490 117.540 ;
        RECT 70.140 117.525 70.370 121.290 ;
        RECT 70.045 117.290 70.370 117.525 ;
        RECT 72.020 117.515 72.250 121.290 ;
        RECT 76.540 119.330 76.890 121.550 ;
        RECT 90.330 121.240 90.560 121.290 ;
        RECT 90.920 121.240 91.150 121.290 ;
        RECT 90.330 121.050 91.150 121.240 ;
        RECT 82.100 119.605 82.330 120.480 ;
        RECT 83.500 119.965 83.730 120.480 ;
        RECT 83.910 119.965 84.910 119.980 ;
        RECT 83.500 119.775 84.910 119.965 ;
        RECT 82.100 119.480 82.525 119.605 ;
        RECT 83.500 119.480 83.730 119.775 ;
        RECT 82.120 119.415 82.525 119.480 ;
        RECT 80.745 119.265 81.035 119.285 ;
        RECT 80.745 119.055 81.305 119.265 ;
        RECT 81.115 118.905 81.305 119.055 ;
        RECT 82.335 118.905 82.525 119.415 ;
        RECT 83.910 118.980 84.910 119.775 ;
        RECT 83.910 118.905 84.100 118.980 ;
        RECT 81.115 118.715 84.100 118.905 ;
        RECT 71.925 117.290 72.250 117.515 ;
        RECT 90.330 117.540 90.560 121.050 ;
        RECT 90.920 117.540 91.150 121.050 ;
        RECT 90.330 117.290 91.150 117.540 ;
        RECT 92.800 117.525 93.030 121.290 ;
        RECT 92.705 117.290 93.030 117.525 ;
        RECT 94.680 117.515 94.910 121.290 ;
        RECT 99.200 119.330 99.550 121.550 ;
        RECT 112.990 121.240 113.220 121.290 ;
        RECT 113.580 121.240 113.810 121.290 ;
        RECT 112.990 121.050 113.810 121.240 ;
        RECT 104.760 119.605 104.990 120.480 ;
        RECT 106.160 119.965 106.390 120.480 ;
        RECT 106.570 119.965 107.570 119.980 ;
        RECT 106.160 119.775 107.570 119.965 ;
        RECT 104.760 119.480 105.185 119.605 ;
        RECT 106.160 119.480 106.390 119.775 ;
        RECT 104.780 119.415 105.185 119.480 ;
        RECT 103.405 119.265 103.695 119.285 ;
        RECT 103.405 119.055 103.965 119.265 ;
        RECT 103.775 118.905 103.965 119.055 ;
        RECT 104.995 118.905 105.185 119.415 ;
        RECT 106.570 118.980 107.570 119.775 ;
        RECT 106.570 118.905 106.760 118.980 ;
        RECT 103.775 118.715 106.760 118.905 ;
        RECT 94.585 117.290 94.910 117.515 ;
        RECT 112.990 117.540 113.220 121.050 ;
        RECT 113.580 117.540 113.810 121.050 ;
        RECT 112.990 117.290 113.810 117.540 ;
        RECT 115.460 117.525 115.690 121.290 ;
        RECT 115.365 117.290 115.690 117.525 ;
        RECT 117.340 117.515 117.570 121.290 ;
        RECT 121.860 119.330 122.210 121.550 ;
        RECT 117.245 117.290 117.570 117.515 ;
        RECT 67.805 116.110 68.365 117.290 ;
        RECT 70.045 116.110 70.235 117.290 ;
        RECT 71.925 116.110 72.115 117.290 ;
        RECT 90.465 116.110 91.025 117.290 ;
        RECT 92.705 116.110 92.895 117.290 ;
        RECT 94.585 116.110 94.775 117.290 ;
        RECT 113.125 116.110 113.685 117.290 ;
        RECT 115.365 116.110 115.555 117.290 ;
        RECT 117.245 116.110 117.435 117.290 ;
        RECT 67.670 115.870 68.490 116.110 ;
        RECT 70.045 115.870 70.370 116.110 ;
        RECT 67.670 112.650 67.900 115.870 ;
        RECT 68.260 112.650 68.490 115.870 ;
        RECT 70.140 112.700 70.370 115.870 ;
        RECT 71.925 115.855 72.250 116.110 ;
        RECT 72.020 112.700 72.250 115.855 ;
        RECT 90.330 115.870 91.150 116.110 ;
        RECT 92.705 115.870 93.030 116.110 ;
        RECT 67.670 112.110 68.490 112.650 ;
        RECT 70.050 112.100 70.650 112.700 ;
        RECT 71.940 112.100 72.540 112.700 ;
        RECT 90.330 112.650 90.560 115.870 ;
        RECT 90.920 112.650 91.150 115.870 ;
        RECT 92.800 112.700 93.030 115.870 ;
        RECT 94.585 115.855 94.910 116.110 ;
        RECT 94.680 112.700 94.910 115.855 ;
        RECT 112.990 115.870 113.810 116.110 ;
        RECT 115.365 115.870 115.690 116.110 ;
        RECT 90.330 112.110 91.150 112.650 ;
        RECT 92.710 112.100 93.310 112.700 ;
        RECT 94.600 112.100 95.200 112.700 ;
        RECT 112.990 112.650 113.220 115.870 ;
        RECT 113.580 112.650 113.810 115.870 ;
        RECT 115.460 112.700 115.690 115.870 ;
        RECT 117.245 115.855 117.570 116.110 ;
        RECT 117.340 112.700 117.570 115.855 ;
        RECT 112.990 112.110 113.810 112.650 ;
        RECT 115.370 112.100 115.970 112.700 ;
        RECT 117.260 112.100 117.860 112.700 ;
        RECT 64.130 111.365 64.460 111.750 ;
        RECT 66.010 111.365 66.340 111.750 ;
        RECT 67.890 111.365 68.220 111.750 ;
        RECT 69.770 111.365 70.100 111.750 ;
        RECT 71.650 111.365 71.980 111.750 ;
        RECT 64.130 111.175 71.980 111.365 ;
        RECT 86.790 111.365 87.120 111.750 ;
        RECT 88.670 111.365 89.000 111.750 ;
        RECT 90.550 111.365 90.880 111.750 ;
        RECT 92.430 111.365 92.760 111.750 ;
        RECT 94.310 111.365 94.640 111.750 ;
        RECT 86.790 111.175 94.640 111.365 ;
        RECT 109.450 111.365 109.780 111.750 ;
        RECT 111.330 111.365 111.660 111.750 ;
        RECT 113.210 111.365 113.540 111.750 ;
        RECT 115.090 111.365 115.420 111.750 ;
        RECT 116.970 111.365 117.300 111.750 ;
        RECT 109.450 111.175 117.300 111.365 ;
        RECT 56.220 107.250 56.570 109.470 ;
        RECT 45.010 103.900 45.240 103.950 ;
        RECT 45.600 103.900 45.830 103.950 ;
        RECT 45.010 103.710 45.830 103.900 ;
        RECT 36.780 102.265 37.010 103.140 ;
        RECT 38.180 102.625 38.410 103.140 ;
        RECT 38.590 102.625 39.590 102.640 ;
        RECT 38.180 102.435 39.590 102.625 ;
        RECT 36.780 102.140 37.205 102.265 ;
        RECT 38.180 102.140 38.410 102.435 ;
        RECT 36.800 102.075 37.205 102.140 ;
        RECT 35.425 101.925 35.715 101.945 ;
        RECT 35.425 101.715 35.985 101.925 ;
        RECT 35.795 101.565 35.985 101.715 ;
        RECT 37.015 101.565 37.205 102.075 ;
        RECT 38.590 101.640 39.590 102.435 ;
        RECT 38.590 101.565 38.780 101.640 ;
        RECT 35.795 101.375 38.780 101.565 ;
        RECT 45.010 100.200 45.240 103.710 ;
        RECT 45.600 100.200 45.830 103.710 ;
        RECT 45.010 99.950 45.830 100.200 ;
        RECT 47.480 100.185 47.710 103.950 ;
        RECT 47.385 99.950 47.710 100.185 ;
        RECT 49.360 100.175 49.590 103.950 ;
        RECT 53.880 101.990 54.230 104.210 ;
        RECT 67.670 103.900 67.900 103.950 ;
        RECT 68.260 103.900 68.490 103.950 ;
        RECT 67.670 103.710 68.490 103.900 ;
        RECT 59.440 102.265 59.670 103.140 ;
        RECT 60.840 102.625 61.070 103.140 ;
        RECT 61.250 102.625 62.250 102.640 ;
        RECT 60.840 102.435 62.250 102.625 ;
        RECT 59.440 102.140 59.865 102.265 ;
        RECT 60.840 102.140 61.070 102.435 ;
        RECT 59.460 102.075 59.865 102.140 ;
        RECT 58.085 101.925 58.375 101.945 ;
        RECT 58.085 101.715 58.645 101.925 ;
        RECT 58.455 101.565 58.645 101.715 ;
        RECT 59.675 101.565 59.865 102.075 ;
        RECT 61.250 101.640 62.250 102.435 ;
        RECT 61.250 101.565 61.440 101.640 ;
        RECT 58.455 101.375 61.440 101.565 ;
        RECT 49.265 99.950 49.590 100.175 ;
        RECT 67.670 100.200 67.900 103.710 ;
        RECT 68.260 100.200 68.490 103.710 ;
        RECT 67.670 99.950 68.490 100.200 ;
        RECT 70.140 100.185 70.370 103.950 ;
        RECT 70.045 99.950 70.370 100.185 ;
        RECT 72.020 100.175 72.250 103.950 ;
        RECT 76.540 101.990 76.890 104.210 ;
        RECT 90.330 103.900 90.560 103.950 ;
        RECT 90.920 103.900 91.150 103.950 ;
        RECT 90.330 103.710 91.150 103.900 ;
        RECT 82.100 102.265 82.330 103.140 ;
        RECT 83.500 102.625 83.730 103.140 ;
        RECT 83.910 102.625 84.910 102.640 ;
        RECT 83.500 102.435 84.910 102.625 ;
        RECT 82.100 102.140 82.525 102.265 ;
        RECT 83.500 102.140 83.730 102.435 ;
        RECT 82.120 102.075 82.525 102.140 ;
        RECT 80.745 101.925 81.035 101.945 ;
        RECT 80.745 101.715 81.305 101.925 ;
        RECT 81.115 101.565 81.305 101.715 ;
        RECT 82.335 101.565 82.525 102.075 ;
        RECT 83.910 101.640 84.910 102.435 ;
        RECT 83.910 101.565 84.100 101.640 ;
        RECT 81.115 101.375 84.100 101.565 ;
        RECT 71.925 99.950 72.250 100.175 ;
        RECT 90.330 100.200 90.560 103.710 ;
        RECT 90.920 100.200 91.150 103.710 ;
        RECT 90.330 99.950 91.150 100.200 ;
        RECT 92.800 100.185 93.030 103.950 ;
        RECT 92.705 99.950 93.030 100.185 ;
        RECT 94.680 100.175 94.910 103.950 ;
        RECT 99.200 101.990 99.550 104.210 ;
        RECT 112.990 103.900 113.220 103.950 ;
        RECT 113.580 103.900 113.810 103.950 ;
        RECT 112.990 103.710 113.810 103.900 ;
        RECT 104.760 102.265 104.990 103.140 ;
        RECT 106.160 102.625 106.390 103.140 ;
        RECT 106.570 102.625 107.570 102.640 ;
        RECT 106.160 102.435 107.570 102.625 ;
        RECT 104.760 102.140 105.185 102.265 ;
        RECT 106.160 102.140 106.390 102.435 ;
        RECT 104.780 102.075 105.185 102.140 ;
        RECT 103.405 101.925 103.695 101.945 ;
        RECT 103.405 101.715 103.965 101.925 ;
        RECT 103.775 101.565 103.965 101.715 ;
        RECT 104.995 101.565 105.185 102.075 ;
        RECT 106.570 101.640 107.570 102.435 ;
        RECT 106.570 101.565 106.760 101.640 ;
        RECT 103.775 101.375 106.760 101.565 ;
        RECT 94.585 99.950 94.910 100.175 ;
        RECT 112.990 100.200 113.220 103.710 ;
        RECT 113.580 100.200 113.810 103.710 ;
        RECT 112.990 99.950 113.810 100.200 ;
        RECT 115.460 100.185 115.690 103.950 ;
        RECT 115.365 99.950 115.690 100.185 ;
        RECT 117.340 100.175 117.570 103.950 ;
        RECT 121.860 101.990 122.210 104.210 ;
        RECT 117.245 99.950 117.570 100.175 ;
        RECT 45.145 98.770 45.705 99.950 ;
        RECT 47.385 98.770 47.575 99.950 ;
        RECT 49.265 98.770 49.455 99.950 ;
        RECT 67.805 98.770 68.365 99.950 ;
        RECT 70.045 98.770 70.235 99.950 ;
        RECT 71.925 98.770 72.115 99.950 ;
        RECT 90.465 98.770 91.025 99.950 ;
        RECT 92.705 98.770 92.895 99.950 ;
        RECT 94.585 98.770 94.775 99.950 ;
        RECT 113.125 98.770 113.685 99.950 ;
        RECT 115.365 98.770 115.555 99.950 ;
        RECT 117.245 98.770 117.435 99.950 ;
        RECT 45.010 98.530 45.830 98.770 ;
        RECT 47.385 98.530 47.710 98.770 ;
        RECT 45.010 95.310 45.240 98.530 ;
        RECT 45.600 95.310 45.830 98.530 ;
        RECT 47.480 95.360 47.710 98.530 ;
        RECT 49.265 98.515 49.590 98.770 ;
        RECT 49.360 95.360 49.590 98.515 ;
        RECT 67.670 98.530 68.490 98.770 ;
        RECT 70.045 98.530 70.370 98.770 ;
        RECT 45.010 94.770 45.830 95.310 ;
        RECT 47.390 94.760 47.990 95.360 ;
        RECT 49.280 94.760 49.880 95.360 ;
        RECT 67.670 95.310 67.900 98.530 ;
        RECT 68.260 95.310 68.490 98.530 ;
        RECT 70.140 95.360 70.370 98.530 ;
        RECT 71.925 98.515 72.250 98.770 ;
        RECT 72.020 95.360 72.250 98.515 ;
        RECT 90.330 98.530 91.150 98.770 ;
        RECT 92.705 98.530 93.030 98.770 ;
        RECT 67.670 94.770 68.490 95.310 ;
        RECT 70.050 94.760 70.650 95.360 ;
        RECT 71.940 94.760 72.540 95.360 ;
        RECT 90.330 95.310 90.560 98.530 ;
        RECT 90.920 95.310 91.150 98.530 ;
        RECT 92.800 95.360 93.030 98.530 ;
        RECT 94.585 98.515 94.910 98.770 ;
        RECT 94.680 95.360 94.910 98.515 ;
        RECT 112.990 98.530 113.810 98.770 ;
        RECT 115.365 98.530 115.690 98.770 ;
        RECT 90.330 94.770 91.150 95.310 ;
        RECT 92.710 94.760 93.310 95.360 ;
        RECT 94.600 94.760 95.200 95.360 ;
        RECT 112.990 95.310 113.220 98.530 ;
        RECT 113.580 95.310 113.810 98.530 ;
        RECT 115.460 95.360 115.690 98.530 ;
        RECT 117.245 98.515 117.570 98.770 ;
        RECT 117.340 95.360 117.570 98.515 ;
        RECT 112.990 94.770 113.810 95.310 ;
        RECT 115.370 94.760 115.970 95.360 ;
        RECT 117.260 94.760 117.860 95.360 ;
        RECT 41.470 94.025 41.800 94.410 ;
        RECT 43.350 94.025 43.680 94.410 ;
        RECT 45.230 94.025 45.560 94.410 ;
        RECT 47.110 94.025 47.440 94.410 ;
        RECT 48.990 94.025 49.320 94.410 ;
        RECT 41.470 93.835 49.320 94.025 ;
        RECT 64.130 94.025 64.460 94.410 ;
        RECT 66.010 94.025 66.340 94.410 ;
        RECT 67.890 94.025 68.220 94.410 ;
        RECT 69.770 94.025 70.100 94.410 ;
        RECT 71.650 94.025 71.980 94.410 ;
        RECT 64.130 93.835 71.980 94.025 ;
        RECT 86.790 94.025 87.120 94.410 ;
        RECT 88.670 94.025 89.000 94.410 ;
        RECT 90.550 94.025 90.880 94.410 ;
        RECT 92.430 94.025 92.760 94.410 ;
        RECT 94.310 94.025 94.640 94.410 ;
        RECT 86.790 93.835 94.640 94.025 ;
        RECT 109.450 94.025 109.780 94.410 ;
        RECT 111.330 94.025 111.660 94.410 ;
        RECT 113.210 94.025 113.540 94.410 ;
        RECT 115.090 94.025 115.420 94.410 ;
        RECT 116.970 94.025 117.300 94.410 ;
        RECT 109.450 93.835 117.300 94.025 ;
        RECT 45.010 86.560 45.240 86.610 ;
        RECT 45.600 86.560 45.830 86.610 ;
        RECT 45.010 86.370 45.830 86.560 ;
        RECT 36.780 84.925 37.010 85.800 ;
        RECT 38.180 85.285 38.410 85.800 ;
        RECT 38.590 85.285 39.590 85.300 ;
        RECT 38.180 85.095 39.590 85.285 ;
        RECT 36.780 84.800 37.205 84.925 ;
        RECT 38.180 84.800 38.410 85.095 ;
        RECT 36.800 84.735 37.205 84.800 ;
        RECT 35.425 84.585 35.715 84.605 ;
        RECT 35.425 84.375 35.985 84.585 ;
        RECT 35.795 84.225 35.985 84.375 ;
        RECT 37.015 84.225 37.205 84.735 ;
        RECT 38.590 84.300 39.590 85.095 ;
        RECT 38.590 84.225 38.780 84.300 ;
        RECT 35.795 84.035 38.780 84.225 ;
        RECT 45.010 82.860 45.240 86.370 ;
        RECT 45.600 82.860 45.830 86.370 ;
        RECT 45.010 82.610 45.830 82.860 ;
        RECT 47.480 82.845 47.710 86.610 ;
        RECT 47.385 82.610 47.710 82.845 ;
        RECT 49.360 82.835 49.590 86.610 ;
        RECT 53.880 84.650 54.230 86.870 ;
        RECT 67.670 86.560 67.900 86.610 ;
        RECT 68.260 86.560 68.490 86.610 ;
        RECT 67.670 86.370 68.490 86.560 ;
        RECT 59.440 84.925 59.670 85.800 ;
        RECT 60.840 85.285 61.070 85.800 ;
        RECT 61.250 85.285 62.250 85.300 ;
        RECT 60.840 85.095 62.250 85.285 ;
        RECT 59.440 84.800 59.865 84.925 ;
        RECT 60.840 84.800 61.070 85.095 ;
        RECT 59.460 84.735 59.865 84.800 ;
        RECT 58.085 84.585 58.375 84.605 ;
        RECT 58.085 84.375 58.645 84.585 ;
        RECT 58.455 84.225 58.645 84.375 ;
        RECT 59.675 84.225 59.865 84.735 ;
        RECT 61.250 84.300 62.250 85.095 ;
        RECT 61.250 84.225 61.440 84.300 ;
        RECT 58.455 84.035 61.440 84.225 ;
        RECT 49.265 82.610 49.590 82.835 ;
        RECT 67.670 82.860 67.900 86.370 ;
        RECT 68.260 82.860 68.490 86.370 ;
        RECT 67.670 82.610 68.490 82.860 ;
        RECT 70.140 82.845 70.370 86.610 ;
        RECT 70.045 82.610 70.370 82.845 ;
        RECT 72.020 82.835 72.250 86.610 ;
        RECT 76.540 84.650 76.890 86.870 ;
        RECT 90.330 86.560 90.560 86.610 ;
        RECT 90.920 86.560 91.150 86.610 ;
        RECT 90.330 86.370 91.150 86.560 ;
        RECT 82.100 84.925 82.330 85.800 ;
        RECT 83.500 85.285 83.730 85.800 ;
        RECT 83.910 85.285 84.910 85.300 ;
        RECT 83.500 85.095 84.910 85.285 ;
        RECT 82.100 84.800 82.525 84.925 ;
        RECT 83.500 84.800 83.730 85.095 ;
        RECT 82.120 84.735 82.525 84.800 ;
        RECT 80.745 84.585 81.035 84.605 ;
        RECT 80.745 84.375 81.305 84.585 ;
        RECT 81.115 84.225 81.305 84.375 ;
        RECT 82.335 84.225 82.525 84.735 ;
        RECT 83.910 84.300 84.910 85.095 ;
        RECT 83.910 84.225 84.100 84.300 ;
        RECT 81.115 84.035 84.100 84.225 ;
        RECT 71.925 82.610 72.250 82.835 ;
        RECT 90.330 82.860 90.560 86.370 ;
        RECT 90.920 82.860 91.150 86.370 ;
        RECT 90.330 82.610 91.150 82.860 ;
        RECT 92.800 82.845 93.030 86.610 ;
        RECT 92.705 82.610 93.030 82.845 ;
        RECT 94.680 82.835 94.910 86.610 ;
        RECT 99.200 84.650 99.550 86.870 ;
        RECT 112.990 86.560 113.220 86.610 ;
        RECT 113.580 86.560 113.810 86.610 ;
        RECT 112.990 86.370 113.810 86.560 ;
        RECT 104.760 84.925 104.990 85.800 ;
        RECT 106.160 85.285 106.390 85.800 ;
        RECT 106.570 85.285 107.570 85.300 ;
        RECT 106.160 85.095 107.570 85.285 ;
        RECT 104.760 84.800 105.185 84.925 ;
        RECT 106.160 84.800 106.390 85.095 ;
        RECT 104.780 84.735 105.185 84.800 ;
        RECT 103.405 84.585 103.695 84.605 ;
        RECT 103.405 84.375 103.965 84.585 ;
        RECT 103.775 84.225 103.965 84.375 ;
        RECT 104.995 84.225 105.185 84.735 ;
        RECT 106.570 84.300 107.570 85.095 ;
        RECT 106.570 84.225 106.760 84.300 ;
        RECT 103.775 84.035 106.760 84.225 ;
        RECT 94.585 82.610 94.910 82.835 ;
        RECT 112.990 82.860 113.220 86.370 ;
        RECT 113.580 82.860 113.810 86.370 ;
        RECT 112.990 82.610 113.810 82.860 ;
        RECT 115.460 82.845 115.690 86.610 ;
        RECT 115.365 82.610 115.690 82.845 ;
        RECT 117.340 82.835 117.570 86.610 ;
        RECT 121.860 84.650 122.210 86.870 ;
        RECT 117.245 82.610 117.570 82.835 ;
        RECT 45.145 81.430 45.705 82.610 ;
        RECT 47.385 81.430 47.575 82.610 ;
        RECT 49.265 81.430 49.455 82.610 ;
        RECT 67.805 81.430 68.365 82.610 ;
        RECT 70.045 81.430 70.235 82.610 ;
        RECT 71.925 81.430 72.115 82.610 ;
        RECT 90.465 81.430 91.025 82.610 ;
        RECT 92.705 81.430 92.895 82.610 ;
        RECT 94.585 81.430 94.775 82.610 ;
        RECT 113.125 81.430 113.685 82.610 ;
        RECT 115.365 81.430 115.555 82.610 ;
        RECT 117.245 81.430 117.435 82.610 ;
        RECT 45.010 81.190 45.830 81.430 ;
        RECT 47.385 81.190 47.710 81.430 ;
        RECT 45.010 77.970 45.240 81.190 ;
        RECT 45.600 77.970 45.830 81.190 ;
        RECT 47.480 78.020 47.710 81.190 ;
        RECT 49.265 81.175 49.590 81.430 ;
        RECT 49.360 78.020 49.590 81.175 ;
        RECT 67.670 81.190 68.490 81.430 ;
        RECT 70.045 81.190 70.370 81.430 ;
        RECT 45.010 77.430 45.830 77.970 ;
        RECT 47.390 77.420 47.990 78.020 ;
        RECT 49.280 77.420 49.880 78.020 ;
        RECT 67.670 77.970 67.900 81.190 ;
        RECT 68.260 77.970 68.490 81.190 ;
        RECT 70.140 78.020 70.370 81.190 ;
        RECT 71.925 81.175 72.250 81.430 ;
        RECT 72.020 78.020 72.250 81.175 ;
        RECT 90.330 81.190 91.150 81.430 ;
        RECT 92.705 81.190 93.030 81.430 ;
        RECT 67.670 77.430 68.490 77.970 ;
        RECT 70.050 77.420 70.650 78.020 ;
        RECT 71.940 77.420 72.540 78.020 ;
        RECT 90.330 77.970 90.560 81.190 ;
        RECT 90.920 77.970 91.150 81.190 ;
        RECT 92.800 78.020 93.030 81.190 ;
        RECT 94.585 81.175 94.910 81.430 ;
        RECT 94.680 78.020 94.910 81.175 ;
        RECT 112.990 81.190 113.810 81.430 ;
        RECT 115.365 81.190 115.690 81.430 ;
        RECT 90.330 77.430 91.150 77.970 ;
        RECT 92.710 77.420 93.310 78.020 ;
        RECT 94.600 77.420 95.200 78.020 ;
        RECT 112.990 77.970 113.220 81.190 ;
        RECT 113.580 77.970 113.810 81.190 ;
        RECT 115.460 78.020 115.690 81.190 ;
        RECT 117.245 81.175 117.570 81.430 ;
        RECT 117.340 78.020 117.570 81.175 ;
        RECT 112.990 77.430 113.810 77.970 ;
        RECT 115.370 77.420 115.970 78.020 ;
        RECT 117.260 77.420 117.860 78.020 ;
        RECT 41.470 76.685 41.800 77.070 ;
        RECT 43.350 76.685 43.680 77.070 ;
        RECT 45.230 76.685 45.560 77.070 ;
        RECT 47.110 76.685 47.440 77.070 ;
        RECT 48.990 76.685 49.320 77.070 ;
        RECT 41.470 76.495 49.320 76.685 ;
        RECT 64.130 76.685 64.460 77.070 ;
        RECT 66.010 76.685 66.340 77.070 ;
        RECT 67.890 76.685 68.220 77.070 ;
        RECT 69.770 76.685 70.100 77.070 ;
        RECT 71.650 76.685 71.980 77.070 ;
        RECT 64.130 76.495 71.980 76.685 ;
        RECT 86.790 76.685 87.120 77.070 ;
        RECT 88.670 76.685 89.000 77.070 ;
        RECT 90.550 76.685 90.880 77.070 ;
        RECT 92.430 76.685 92.760 77.070 ;
        RECT 94.310 76.685 94.640 77.070 ;
        RECT 86.790 76.495 94.640 76.685 ;
        RECT 109.450 76.685 109.780 77.070 ;
        RECT 111.330 76.685 111.660 77.070 ;
        RECT 113.210 76.685 113.540 77.070 ;
        RECT 115.090 76.685 115.420 77.070 ;
        RECT 116.970 76.685 117.300 77.070 ;
        RECT 109.450 76.495 117.300 76.685 ;
        RECT 45.010 69.220 45.240 69.270 ;
        RECT 45.600 69.220 45.830 69.270 ;
        RECT 45.010 69.030 45.830 69.220 ;
        RECT 36.780 67.585 37.010 68.460 ;
        RECT 38.180 67.945 38.410 68.460 ;
        RECT 38.590 67.945 39.590 67.960 ;
        RECT 38.180 67.755 39.590 67.945 ;
        RECT 36.780 67.460 37.205 67.585 ;
        RECT 38.180 67.460 38.410 67.755 ;
        RECT 36.800 67.395 37.205 67.460 ;
        RECT 35.425 67.245 35.715 67.265 ;
        RECT 35.425 67.035 35.985 67.245 ;
        RECT 35.795 66.885 35.985 67.035 ;
        RECT 37.015 66.885 37.205 67.395 ;
        RECT 38.590 66.960 39.590 67.755 ;
        RECT 38.590 66.885 38.780 66.960 ;
        RECT 35.795 66.695 38.780 66.885 ;
        RECT 45.010 65.520 45.240 69.030 ;
        RECT 45.600 65.520 45.830 69.030 ;
        RECT 45.010 65.270 45.830 65.520 ;
        RECT 47.480 65.505 47.710 69.270 ;
        RECT 47.385 65.270 47.710 65.505 ;
        RECT 49.360 65.495 49.590 69.270 ;
        RECT 53.880 67.310 54.230 69.530 ;
        RECT 67.670 69.220 67.900 69.270 ;
        RECT 68.260 69.220 68.490 69.270 ;
        RECT 67.670 69.030 68.490 69.220 ;
        RECT 59.440 67.585 59.670 68.460 ;
        RECT 60.840 67.945 61.070 68.460 ;
        RECT 61.250 67.945 62.250 67.960 ;
        RECT 60.840 67.755 62.250 67.945 ;
        RECT 59.440 67.460 59.865 67.585 ;
        RECT 60.840 67.460 61.070 67.755 ;
        RECT 59.460 67.395 59.865 67.460 ;
        RECT 58.085 67.245 58.375 67.265 ;
        RECT 58.085 67.035 58.645 67.245 ;
        RECT 58.455 66.885 58.645 67.035 ;
        RECT 59.675 66.885 59.865 67.395 ;
        RECT 61.250 66.960 62.250 67.755 ;
        RECT 61.250 66.885 61.440 66.960 ;
        RECT 58.455 66.695 61.440 66.885 ;
        RECT 49.265 65.270 49.590 65.495 ;
        RECT 67.670 65.520 67.900 69.030 ;
        RECT 68.260 65.520 68.490 69.030 ;
        RECT 67.670 65.270 68.490 65.520 ;
        RECT 70.140 65.505 70.370 69.270 ;
        RECT 70.045 65.270 70.370 65.505 ;
        RECT 72.020 65.495 72.250 69.270 ;
        RECT 76.540 67.310 76.890 69.530 ;
        RECT 90.330 69.220 90.560 69.270 ;
        RECT 90.920 69.220 91.150 69.270 ;
        RECT 90.330 69.030 91.150 69.220 ;
        RECT 82.100 67.585 82.330 68.460 ;
        RECT 83.500 67.945 83.730 68.460 ;
        RECT 83.910 67.945 84.910 67.960 ;
        RECT 83.500 67.755 84.910 67.945 ;
        RECT 82.100 67.460 82.525 67.585 ;
        RECT 83.500 67.460 83.730 67.755 ;
        RECT 82.120 67.395 82.525 67.460 ;
        RECT 80.745 67.245 81.035 67.265 ;
        RECT 80.745 67.035 81.305 67.245 ;
        RECT 81.115 66.885 81.305 67.035 ;
        RECT 82.335 66.885 82.525 67.395 ;
        RECT 83.910 66.960 84.910 67.755 ;
        RECT 83.910 66.885 84.100 66.960 ;
        RECT 81.115 66.695 84.100 66.885 ;
        RECT 71.925 65.270 72.250 65.495 ;
        RECT 90.330 65.520 90.560 69.030 ;
        RECT 90.920 65.520 91.150 69.030 ;
        RECT 90.330 65.270 91.150 65.520 ;
        RECT 92.800 65.505 93.030 69.270 ;
        RECT 92.705 65.270 93.030 65.505 ;
        RECT 94.680 65.495 94.910 69.270 ;
        RECT 99.200 67.310 99.550 69.530 ;
        RECT 112.990 69.220 113.220 69.270 ;
        RECT 113.580 69.220 113.810 69.270 ;
        RECT 112.990 69.030 113.810 69.220 ;
        RECT 104.760 67.585 104.990 68.460 ;
        RECT 106.160 67.945 106.390 68.460 ;
        RECT 106.570 67.945 107.570 67.960 ;
        RECT 106.160 67.755 107.570 67.945 ;
        RECT 104.760 67.460 105.185 67.585 ;
        RECT 106.160 67.460 106.390 67.755 ;
        RECT 104.780 67.395 105.185 67.460 ;
        RECT 103.405 67.245 103.695 67.265 ;
        RECT 103.405 67.035 103.965 67.245 ;
        RECT 103.775 66.885 103.965 67.035 ;
        RECT 104.995 66.885 105.185 67.395 ;
        RECT 106.570 66.960 107.570 67.755 ;
        RECT 106.570 66.885 106.760 66.960 ;
        RECT 103.775 66.695 106.760 66.885 ;
        RECT 94.585 65.270 94.910 65.495 ;
        RECT 112.990 65.520 113.220 69.030 ;
        RECT 113.580 65.520 113.810 69.030 ;
        RECT 112.990 65.270 113.810 65.520 ;
        RECT 115.460 65.505 115.690 69.270 ;
        RECT 115.365 65.270 115.690 65.505 ;
        RECT 117.340 65.495 117.570 69.270 ;
        RECT 121.860 67.310 122.210 69.530 ;
        RECT 117.245 65.270 117.570 65.495 ;
        RECT 45.145 64.090 45.705 65.270 ;
        RECT 47.385 64.090 47.575 65.270 ;
        RECT 49.265 64.090 49.455 65.270 ;
        RECT 67.805 64.090 68.365 65.270 ;
        RECT 70.045 64.090 70.235 65.270 ;
        RECT 71.925 64.090 72.115 65.270 ;
        RECT 90.465 64.090 91.025 65.270 ;
        RECT 92.705 64.090 92.895 65.270 ;
        RECT 94.585 64.090 94.775 65.270 ;
        RECT 113.125 64.090 113.685 65.270 ;
        RECT 115.365 64.090 115.555 65.270 ;
        RECT 117.245 64.090 117.435 65.270 ;
        RECT 45.010 63.850 45.830 64.090 ;
        RECT 47.385 63.850 47.710 64.090 ;
        RECT 45.010 60.630 45.240 63.850 ;
        RECT 45.600 60.630 45.830 63.850 ;
        RECT 47.480 60.680 47.710 63.850 ;
        RECT 49.265 63.835 49.590 64.090 ;
        RECT 49.360 60.680 49.590 63.835 ;
        RECT 67.670 63.850 68.490 64.090 ;
        RECT 70.045 63.850 70.370 64.090 ;
        RECT 45.010 60.090 45.830 60.630 ;
        RECT 47.390 60.080 47.990 60.680 ;
        RECT 49.280 60.080 49.880 60.680 ;
        RECT 67.670 60.630 67.900 63.850 ;
        RECT 68.260 60.630 68.490 63.850 ;
        RECT 70.140 60.680 70.370 63.850 ;
        RECT 71.925 63.835 72.250 64.090 ;
        RECT 72.020 60.680 72.250 63.835 ;
        RECT 90.330 63.850 91.150 64.090 ;
        RECT 92.705 63.850 93.030 64.090 ;
        RECT 67.670 60.090 68.490 60.630 ;
        RECT 70.050 60.080 70.650 60.680 ;
        RECT 71.940 60.080 72.540 60.680 ;
        RECT 90.330 60.630 90.560 63.850 ;
        RECT 90.920 60.630 91.150 63.850 ;
        RECT 92.800 60.680 93.030 63.850 ;
        RECT 94.585 63.835 94.910 64.090 ;
        RECT 94.680 60.680 94.910 63.835 ;
        RECT 112.990 63.850 113.810 64.090 ;
        RECT 115.365 63.850 115.690 64.090 ;
        RECT 90.330 60.090 91.150 60.630 ;
        RECT 92.710 60.080 93.310 60.680 ;
        RECT 94.600 60.080 95.200 60.680 ;
        RECT 112.990 60.630 113.220 63.850 ;
        RECT 113.580 60.630 113.810 63.850 ;
        RECT 115.460 60.680 115.690 63.850 ;
        RECT 117.245 63.835 117.570 64.090 ;
        RECT 117.340 60.680 117.570 63.835 ;
        RECT 112.990 60.090 113.810 60.630 ;
        RECT 115.370 60.080 115.970 60.680 ;
        RECT 117.260 60.080 117.860 60.680 ;
        RECT 41.470 59.345 41.800 59.730 ;
        RECT 43.350 59.345 43.680 59.730 ;
        RECT 45.230 59.345 45.560 59.730 ;
        RECT 47.110 59.345 47.440 59.730 ;
        RECT 48.990 59.345 49.320 59.730 ;
        RECT 41.470 59.155 49.320 59.345 ;
        RECT 64.130 59.345 64.460 59.730 ;
        RECT 66.010 59.345 66.340 59.730 ;
        RECT 67.890 59.345 68.220 59.730 ;
        RECT 69.770 59.345 70.100 59.730 ;
        RECT 71.650 59.345 71.980 59.730 ;
        RECT 64.130 59.155 71.980 59.345 ;
        RECT 86.790 59.345 87.120 59.730 ;
        RECT 88.670 59.345 89.000 59.730 ;
        RECT 90.550 59.345 90.880 59.730 ;
        RECT 92.430 59.345 92.760 59.730 ;
        RECT 94.310 59.345 94.640 59.730 ;
        RECT 86.790 59.155 94.640 59.345 ;
        RECT 109.450 59.345 109.780 59.730 ;
        RECT 111.330 59.345 111.660 59.730 ;
        RECT 113.210 59.345 113.540 59.730 ;
        RECT 115.090 59.345 115.420 59.730 ;
        RECT 116.970 59.345 117.300 59.730 ;
        RECT 109.450 59.155 117.300 59.345 ;
        RECT 45.010 51.220 45.240 51.270 ;
        RECT 45.600 51.220 45.830 51.270 ;
        RECT 45.010 51.030 45.830 51.220 ;
        RECT 45.010 47.520 45.240 51.030 ;
        RECT 45.600 47.520 45.830 51.030 ;
        RECT 45.010 47.270 45.830 47.520 ;
        RECT 47.480 47.505 47.710 51.270 ;
        RECT 47.385 47.270 47.710 47.505 ;
        RECT 49.360 47.495 49.590 51.270 ;
        RECT 53.880 49.310 54.230 51.530 ;
        RECT 67.670 51.220 67.900 51.270 ;
        RECT 68.260 51.220 68.490 51.270 ;
        RECT 67.670 51.030 68.490 51.220 ;
        RECT 49.265 47.270 49.590 47.495 ;
        RECT 67.670 47.520 67.900 51.030 ;
        RECT 68.260 47.520 68.490 51.030 ;
        RECT 67.670 47.270 68.490 47.520 ;
        RECT 70.140 47.505 70.370 51.270 ;
        RECT 70.045 47.270 70.370 47.505 ;
        RECT 72.020 47.495 72.250 51.270 ;
        RECT 76.540 49.310 76.890 51.530 ;
        RECT 90.330 51.220 90.560 51.270 ;
        RECT 90.920 51.220 91.150 51.270 ;
        RECT 90.330 51.030 91.150 51.220 ;
        RECT 71.925 47.270 72.250 47.495 ;
        RECT 90.330 47.520 90.560 51.030 ;
        RECT 90.920 47.520 91.150 51.030 ;
        RECT 90.330 47.270 91.150 47.520 ;
        RECT 92.800 47.505 93.030 51.270 ;
        RECT 92.705 47.270 93.030 47.505 ;
        RECT 94.680 47.495 94.910 51.270 ;
        RECT 99.200 49.310 99.550 51.530 ;
        RECT 112.990 51.220 113.220 51.270 ;
        RECT 113.580 51.220 113.810 51.270 ;
        RECT 112.990 51.030 113.810 51.220 ;
        RECT 94.585 47.270 94.910 47.495 ;
        RECT 112.990 47.520 113.220 51.030 ;
        RECT 113.580 47.520 113.810 51.030 ;
        RECT 112.990 47.270 113.810 47.520 ;
        RECT 115.460 47.505 115.690 51.270 ;
        RECT 115.365 47.270 115.690 47.505 ;
        RECT 117.340 47.495 117.570 51.270 ;
        RECT 121.860 49.310 122.210 51.530 ;
        RECT 117.245 47.270 117.570 47.495 ;
        RECT 45.145 46.090 45.705 47.270 ;
        RECT 47.385 46.090 47.575 47.270 ;
        RECT 49.265 46.090 49.455 47.270 ;
        RECT 67.805 46.090 68.365 47.270 ;
        RECT 70.045 46.090 70.235 47.270 ;
        RECT 71.925 46.090 72.115 47.270 ;
        RECT 90.465 46.090 91.025 47.270 ;
        RECT 92.705 46.090 92.895 47.270 ;
        RECT 94.585 46.090 94.775 47.270 ;
        RECT 113.125 46.090 113.685 47.270 ;
        RECT 115.365 46.090 115.555 47.270 ;
        RECT 117.245 46.090 117.435 47.270 ;
        RECT 45.010 45.850 45.830 46.090 ;
        RECT 47.385 45.850 47.710 46.090 ;
        RECT 45.010 42.630 45.240 45.850 ;
        RECT 45.600 42.630 45.830 45.850 ;
        RECT 47.480 42.680 47.710 45.850 ;
        RECT 49.265 45.835 49.590 46.090 ;
        RECT 49.360 42.680 49.590 45.835 ;
        RECT 67.670 45.850 68.490 46.090 ;
        RECT 70.045 45.850 70.370 46.090 ;
        RECT 45.010 42.090 45.830 42.630 ;
        RECT 47.390 42.080 47.990 42.680 ;
        RECT 49.280 42.080 49.880 42.680 ;
        RECT 67.670 42.630 67.900 45.850 ;
        RECT 68.260 42.630 68.490 45.850 ;
        RECT 70.140 42.680 70.370 45.850 ;
        RECT 71.925 45.835 72.250 46.090 ;
        RECT 72.020 42.680 72.250 45.835 ;
        RECT 90.330 45.850 91.150 46.090 ;
        RECT 92.705 45.850 93.030 46.090 ;
        RECT 67.670 42.090 68.490 42.630 ;
        RECT 70.050 42.080 70.650 42.680 ;
        RECT 71.940 42.080 72.540 42.680 ;
        RECT 90.330 42.630 90.560 45.850 ;
        RECT 90.920 42.630 91.150 45.850 ;
        RECT 92.800 42.680 93.030 45.850 ;
        RECT 94.585 45.835 94.910 46.090 ;
        RECT 94.680 42.680 94.910 45.835 ;
        RECT 112.990 45.850 113.810 46.090 ;
        RECT 115.365 45.850 115.690 46.090 ;
        RECT 90.330 42.090 91.150 42.630 ;
        RECT 92.710 42.080 93.310 42.680 ;
        RECT 94.600 42.080 95.200 42.680 ;
        RECT 112.990 42.630 113.220 45.850 ;
        RECT 113.580 42.630 113.810 45.850 ;
        RECT 115.460 42.680 115.690 45.850 ;
        RECT 117.245 45.835 117.570 46.090 ;
        RECT 117.340 42.680 117.570 45.835 ;
        RECT 112.990 42.090 113.810 42.630 ;
        RECT 115.370 42.080 115.970 42.680 ;
        RECT 117.260 42.080 117.860 42.680 ;
        RECT 41.470 41.345 41.800 41.730 ;
        RECT 43.350 41.345 43.680 41.730 ;
        RECT 45.230 41.345 45.560 41.730 ;
        RECT 47.110 41.345 47.440 41.730 ;
        RECT 48.990 41.345 49.320 41.730 ;
        RECT 41.470 41.155 49.320 41.345 ;
        RECT 64.130 41.345 64.460 41.730 ;
        RECT 66.010 41.345 66.340 41.730 ;
        RECT 67.890 41.345 68.220 41.730 ;
        RECT 69.770 41.345 70.100 41.730 ;
        RECT 71.650 41.345 71.980 41.730 ;
        RECT 64.130 41.155 71.980 41.345 ;
        RECT 86.790 41.345 87.120 41.730 ;
        RECT 88.670 41.345 89.000 41.730 ;
        RECT 90.550 41.345 90.880 41.730 ;
        RECT 92.430 41.345 92.760 41.730 ;
        RECT 94.310 41.345 94.640 41.730 ;
        RECT 86.790 41.155 94.640 41.345 ;
        RECT 109.450 41.345 109.780 41.730 ;
        RECT 111.330 41.345 111.660 41.730 ;
        RECT 113.210 41.345 113.540 41.730 ;
        RECT 115.090 41.345 115.420 41.730 ;
        RECT 116.970 41.345 117.300 41.730 ;
        RECT 109.450 41.155 117.300 41.345 ;
      LAYER via ;
        RECT 50.265 186.460 50.525 186.720 ;
        RECT 50.585 186.460 50.845 186.720 ;
        RECT 50.905 186.460 51.165 186.720 ;
        RECT 51.225 186.460 51.485 186.720 ;
        RECT 51.545 186.460 51.805 186.720 ;
        RECT 68.775 186.460 69.035 186.720 ;
        RECT 69.095 186.460 69.355 186.720 ;
        RECT 69.415 186.460 69.675 186.720 ;
        RECT 69.735 186.460 69.995 186.720 ;
        RECT 70.055 186.460 70.315 186.720 ;
        RECT 87.285 186.460 87.545 186.720 ;
        RECT 87.605 186.460 87.865 186.720 ;
        RECT 87.925 186.460 88.185 186.720 ;
        RECT 88.245 186.460 88.505 186.720 ;
        RECT 88.565 186.460 88.825 186.720 ;
        RECT 105.795 186.460 106.055 186.720 ;
        RECT 106.115 186.460 106.375 186.720 ;
        RECT 106.435 186.460 106.695 186.720 ;
        RECT 106.755 186.460 107.015 186.720 ;
        RECT 107.075 186.460 107.335 186.720 ;
        RECT 50.265 181.020 50.525 181.280 ;
        RECT 50.585 181.020 50.845 181.280 ;
        RECT 50.905 181.020 51.165 181.280 ;
        RECT 51.225 181.020 51.485 181.280 ;
        RECT 51.545 181.020 51.805 181.280 ;
        RECT 68.775 181.020 69.035 181.280 ;
        RECT 69.095 181.020 69.355 181.280 ;
        RECT 69.415 181.020 69.675 181.280 ;
        RECT 69.735 181.020 69.995 181.280 ;
        RECT 70.055 181.020 70.315 181.280 ;
        RECT 87.285 181.020 87.545 181.280 ;
        RECT 87.605 181.020 87.865 181.280 ;
        RECT 87.925 181.020 88.185 181.280 ;
        RECT 88.245 181.020 88.505 181.280 ;
        RECT 88.565 181.020 88.825 181.280 ;
        RECT 105.795 181.020 106.055 181.280 ;
        RECT 106.115 181.020 106.375 181.280 ;
        RECT 106.435 181.020 106.695 181.280 ;
        RECT 106.755 181.020 107.015 181.280 ;
        RECT 107.075 181.020 107.335 181.280 ;
        RECT 50.265 175.580 50.525 175.840 ;
        RECT 50.585 175.580 50.845 175.840 ;
        RECT 50.905 175.580 51.165 175.840 ;
        RECT 51.225 175.580 51.485 175.840 ;
        RECT 51.545 175.580 51.805 175.840 ;
        RECT 68.775 175.580 69.035 175.840 ;
        RECT 69.095 175.580 69.355 175.840 ;
        RECT 69.415 175.580 69.675 175.840 ;
        RECT 69.735 175.580 69.995 175.840 ;
        RECT 70.055 175.580 70.315 175.840 ;
        RECT 87.285 175.580 87.545 175.840 ;
        RECT 87.605 175.580 87.865 175.840 ;
        RECT 87.925 175.580 88.185 175.840 ;
        RECT 88.245 175.580 88.505 175.840 ;
        RECT 88.565 175.580 88.825 175.840 ;
        RECT 105.795 175.580 106.055 175.840 ;
        RECT 106.115 175.580 106.375 175.840 ;
        RECT 106.435 175.580 106.695 175.840 ;
        RECT 106.755 175.580 107.015 175.840 ;
        RECT 107.075 175.580 107.335 175.840 ;
        RECT 50.265 170.140 50.525 170.400 ;
        RECT 50.585 170.140 50.845 170.400 ;
        RECT 50.905 170.140 51.165 170.400 ;
        RECT 51.225 170.140 51.485 170.400 ;
        RECT 51.545 170.140 51.805 170.400 ;
        RECT 68.775 170.140 69.035 170.400 ;
        RECT 69.095 170.140 69.355 170.400 ;
        RECT 69.415 170.140 69.675 170.400 ;
        RECT 69.735 170.140 69.995 170.400 ;
        RECT 70.055 170.140 70.315 170.400 ;
        RECT 87.285 170.140 87.545 170.400 ;
        RECT 87.605 170.140 87.865 170.400 ;
        RECT 87.925 170.140 88.185 170.400 ;
        RECT 88.245 170.140 88.505 170.400 ;
        RECT 88.565 170.140 88.825 170.400 ;
        RECT 105.795 170.140 106.055 170.400 ;
        RECT 106.115 170.140 106.375 170.400 ;
        RECT 106.435 170.140 106.695 170.400 ;
        RECT 106.755 170.140 107.015 170.400 ;
        RECT 107.075 170.140 107.335 170.400 ;
        RECT 50.265 164.700 50.525 164.960 ;
        RECT 50.585 164.700 50.845 164.960 ;
        RECT 50.905 164.700 51.165 164.960 ;
        RECT 51.225 164.700 51.485 164.960 ;
        RECT 51.545 164.700 51.805 164.960 ;
        RECT 68.775 164.700 69.035 164.960 ;
        RECT 69.095 164.700 69.355 164.960 ;
        RECT 69.415 164.700 69.675 164.960 ;
        RECT 69.735 164.700 69.995 164.960 ;
        RECT 70.055 164.700 70.315 164.960 ;
        RECT 87.285 164.700 87.545 164.960 ;
        RECT 87.605 164.700 87.865 164.960 ;
        RECT 87.925 164.700 88.185 164.960 ;
        RECT 88.245 164.700 88.505 164.960 ;
        RECT 88.565 164.700 88.825 164.960 ;
        RECT 105.795 164.700 106.055 164.960 ;
        RECT 106.115 164.700 106.375 164.960 ;
        RECT 106.435 164.700 106.695 164.960 ;
        RECT 106.755 164.700 107.015 164.960 ;
        RECT 107.075 164.700 107.335 164.960 ;
        RECT 50.265 159.260 50.525 159.520 ;
        RECT 50.585 159.260 50.845 159.520 ;
        RECT 50.905 159.260 51.165 159.520 ;
        RECT 51.225 159.260 51.485 159.520 ;
        RECT 51.545 159.260 51.805 159.520 ;
        RECT 68.775 159.260 69.035 159.520 ;
        RECT 69.095 159.260 69.355 159.520 ;
        RECT 69.415 159.260 69.675 159.520 ;
        RECT 69.735 159.260 69.995 159.520 ;
        RECT 70.055 159.260 70.315 159.520 ;
        RECT 87.285 159.260 87.545 159.520 ;
        RECT 87.605 159.260 87.865 159.520 ;
        RECT 87.925 159.260 88.185 159.520 ;
        RECT 88.245 159.260 88.505 159.520 ;
        RECT 88.565 159.260 88.825 159.520 ;
        RECT 105.795 159.260 106.055 159.520 ;
        RECT 106.115 159.260 106.375 159.520 ;
        RECT 106.435 159.260 106.695 159.520 ;
        RECT 106.755 159.260 107.015 159.520 ;
        RECT 107.075 159.260 107.335 159.520 ;
        RECT 61.290 119.020 62.210 119.940 ;
        RECT 76.540 119.360 76.890 121.520 ;
        RECT 83.950 119.020 84.870 119.940 ;
        RECT 99.200 119.360 99.550 121.520 ;
        RECT 106.610 119.020 107.530 119.940 ;
        RECT 121.860 119.360 122.210 121.520 ;
        RECT 67.700 112.140 68.450 112.620 ;
        RECT 70.080 112.130 70.620 112.670 ;
        RECT 71.970 112.130 72.510 112.670 ;
        RECT 90.360 112.140 91.110 112.620 ;
        RECT 92.740 112.130 93.280 112.670 ;
        RECT 94.630 112.130 95.170 112.670 ;
        RECT 113.020 112.140 113.770 112.620 ;
        RECT 115.400 112.130 115.940 112.670 ;
        RECT 117.290 112.130 117.830 112.670 ;
        RECT 71.685 111.450 71.945 111.710 ;
        RECT 94.345 111.450 94.605 111.710 ;
        RECT 117.005 111.450 117.265 111.710 ;
        RECT 56.220 107.280 56.570 109.440 ;
        RECT 38.630 101.680 39.550 102.600 ;
        RECT 53.880 102.020 54.230 104.180 ;
        RECT 61.290 101.680 62.210 102.600 ;
        RECT 76.540 102.020 76.890 104.180 ;
        RECT 83.950 101.680 84.870 102.600 ;
        RECT 99.200 102.020 99.550 104.180 ;
        RECT 106.610 101.680 107.530 102.600 ;
        RECT 121.860 102.020 122.210 104.180 ;
        RECT 45.040 94.800 45.790 95.280 ;
        RECT 47.420 94.790 47.960 95.330 ;
        RECT 49.310 94.790 49.850 95.330 ;
        RECT 67.700 94.800 68.450 95.280 ;
        RECT 70.080 94.790 70.620 95.330 ;
        RECT 71.970 94.790 72.510 95.330 ;
        RECT 90.360 94.800 91.110 95.280 ;
        RECT 92.740 94.790 93.280 95.330 ;
        RECT 94.630 94.790 95.170 95.330 ;
        RECT 113.020 94.800 113.770 95.280 ;
        RECT 115.400 94.790 115.940 95.330 ;
        RECT 117.290 94.790 117.830 95.330 ;
        RECT 49.025 94.110 49.285 94.370 ;
        RECT 71.685 94.110 71.945 94.370 ;
        RECT 94.345 94.110 94.605 94.370 ;
        RECT 117.005 94.110 117.265 94.370 ;
        RECT 38.630 84.340 39.550 85.260 ;
        RECT 53.880 84.680 54.230 86.840 ;
        RECT 61.290 84.340 62.210 85.260 ;
        RECT 76.540 84.680 76.890 86.840 ;
        RECT 83.950 84.340 84.870 85.260 ;
        RECT 99.200 84.680 99.550 86.840 ;
        RECT 106.610 84.340 107.530 85.260 ;
        RECT 121.860 84.680 122.210 86.840 ;
        RECT 45.040 77.460 45.790 77.940 ;
        RECT 47.420 77.450 47.960 77.990 ;
        RECT 49.310 77.450 49.850 77.990 ;
        RECT 67.700 77.460 68.450 77.940 ;
        RECT 70.080 77.450 70.620 77.990 ;
        RECT 71.970 77.450 72.510 77.990 ;
        RECT 90.360 77.460 91.110 77.940 ;
        RECT 92.740 77.450 93.280 77.990 ;
        RECT 94.630 77.450 95.170 77.990 ;
        RECT 113.020 77.460 113.770 77.940 ;
        RECT 115.400 77.450 115.940 77.990 ;
        RECT 117.290 77.450 117.830 77.990 ;
        RECT 49.025 76.770 49.285 77.030 ;
        RECT 71.685 76.770 71.945 77.030 ;
        RECT 94.345 76.770 94.605 77.030 ;
        RECT 117.005 76.770 117.265 77.030 ;
        RECT 38.630 67.000 39.550 67.920 ;
        RECT 53.880 67.340 54.230 69.500 ;
        RECT 61.290 67.000 62.210 67.920 ;
        RECT 76.540 67.340 76.890 69.500 ;
        RECT 83.950 67.000 84.870 67.920 ;
        RECT 99.200 67.340 99.550 69.500 ;
        RECT 106.610 67.000 107.530 67.920 ;
        RECT 121.860 67.340 122.210 69.500 ;
        RECT 45.040 60.120 45.790 60.600 ;
        RECT 47.420 60.110 47.960 60.650 ;
        RECT 49.310 60.110 49.850 60.650 ;
        RECT 67.700 60.120 68.450 60.600 ;
        RECT 70.080 60.110 70.620 60.650 ;
        RECT 71.970 60.110 72.510 60.650 ;
        RECT 90.360 60.120 91.110 60.600 ;
        RECT 92.740 60.110 93.280 60.650 ;
        RECT 94.630 60.110 95.170 60.650 ;
        RECT 113.020 60.120 113.770 60.600 ;
        RECT 115.400 60.110 115.940 60.650 ;
        RECT 117.290 60.110 117.830 60.650 ;
        RECT 49.025 59.430 49.285 59.690 ;
        RECT 71.685 59.430 71.945 59.690 ;
        RECT 94.345 59.430 94.605 59.690 ;
        RECT 117.005 59.430 117.265 59.690 ;
        RECT 53.880 49.340 54.230 51.500 ;
        RECT 76.540 49.340 76.890 51.500 ;
        RECT 99.200 49.340 99.550 51.500 ;
        RECT 121.860 49.340 122.210 51.500 ;
        RECT 45.040 42.120 45.790 42.600 ;
        RECT 47.420 42.110 47.960 42.650 ;
        RECT 49.310 42.110 49.850 42.650 ;
        RECT 67.700 42.120 68.450 42.600 ;
        RECT 70.080 42.110 70.620 42.650 ;
        RECT 71.970 42.110 72.510 42.650 ;
        RECT 90.360 42.120 91.110 42.600 ;
        RECT 92.740 42.110 93.280 42.650 ;
        RECT 94.630 42.110 95.170 42.650 ;
        RECT 113.020 42.120 113.770 42.600 ;
        RECT 115.400 42.110 115.940 42.650 ;
        RECT 117.290 42.110 117.830 42.650 ;
        RECT 49.025 41.430 49.285 41.690 ;
        RECT 71.685 41.430 71.945 41.690 ;
        RECT 94.345 41.430 94.605 41.690 ;
        RECT 117.005 41.430 117.265 41.690 ;
      LAYER met2 ;
        RECT 50.265 186.405 51.805 186.775 ;
        RECT 68.775 186.405 70.315 186.775 ;
        RECT 87.285 186.405 88.825 186.775 ;
        RECT 105.795 186.405 107.335 186.775 ;
        RECT 50.265 180.965 51.805 181.335 ;
        RECT 68.775 180.965 70.315 181.335 ;
        RECT 87.285 180.965 88.825 181.335 ;
        RECT 105.795 180.965 107.335 181.335 ;
        RECT 50.265 175.525 51.805 175.895 ;
        RECT 68.775 175.525 70.315 175.895 ;
        RECT 87.285 175.525 88.825 175.895 ;
        RECT 105.795 175.525 107.335 175.895 ;
        RECT 50.265 170.085 51.805 170.455 ;
        RECT 68.775 170.085 70.315 170.455 ;
        RECT 87.285 170.085 88.825 170.455 ;
        RECT 105.795 170.085 107.335 170.455 ;
        RECT 50.265 164.645 51.805 165.015 ;
        RECT 68.775 164.645 70.315 165.015 ;
        RECT 87.285 164.645 88.825 165.015 ;
        RECT 105.795 164.645 107.335 165.015 ;
        RECT 50.265 159.205 51.805 159.575 ;
        RECT 68.775 159.205 70.315 159.575 ;
        RECT 87.285 159.205 88.825 159.575 ;
        RECT 105.795 159.205 107.335 159.575 ;
        RECT 75.890 121.870 76.890 122.870 ;
        RECT 98.550 121.870 99.550 122.870 ;
        RECT 121.210 121.870 122.210 122.870 ;
        RECT 76.590 121.550 76.840 121.870 ;
        RECT 99.250 121.550 99.500 121.870 ;
        RECT 121.910 121.550 122.160 121.870 ;
        RECT 61.250 119.270 62.250 119.980 ;
        RECT 76.540 119.330 76.890 121.550 ;
        RECT 61.250 119.030 62.720 119.270 ;
        RECT 61.250 118.980 62.250 119.030 ;
        RECT 32.920 46.125 33.920 117.245 ;
        RECT 62.480 112.500 62.720 119.030 ;
        RECT 67.590 112.500 68.590 113.110 ;
        RECT 69.650 112.500 70.650 113.100 ;
        RECT 71.540 112.500 72.540 113.100 ;
        RECT 76.600 112.500 76.840 119.330 ;
        RECT 83.910 119.270 84.910 119.980 ;
        RECT 99.200 119.330 99.550 121.550 ;
        RECT 83.910 119.030 85.380 119.270 ;
        RECT 83.910 118.980 84.910 119.030 ;
        RECT 62.480 112.260 76.840 112.500 ;
        RECT 85.140 112.500 85.380 119.030 ;
        RECT 90.250 112.500 91.250 113.110 ;
        RECT 92.310 112.500 93.310 113.100 ;
        RECT 94.200 112.500 95.200 113.100 ;
        RECT 99.260 112.500 99.500 119.330 ;
        RECT 106.570 119.270 107.570 119.980 ;
        RECT 121.860 119.330 122.210 121.550 ;
        RECT 106.570 119.030 108.040 119.270 ;
        RECT 106.570 118.980 107.570 119.030 ;
        RECT 85.140 112.260 99.500 112.500 ;
        RECT 107.800 112.500 108.040 119.030 ;
        RECT 112.910 112.500 113.910 113.110 ;
        RECT 114.970 112.500 115.970 113.100 ;
        RECT 116.860 112.500 117.860 113.100 ;
        RECT 121.920 112.500 122.160 119.330 ;
        RECT 125.830 117.165 126.830 117.190 ;
        RECT 125.810 116.215 126.850 117.165 ;
        RECT 107.800 112.260 122.160 112.500 ;
        RECT 67.590 112.110 68.590 112.260 ;
        RECT 69.650 112.100 70.650 112.260 ;
        RECT 71.540 112.100 72.540 112.260 ;
        RECT 90.250 112.110 91.250 112.260 ;
        RECT 92.310 112.100 93.310 112.260 ;
        RECT 94.200 112.100 95.200 112.260 ;
        RECT 112.910 112.110 113.910 112.260 ;
        RECT 114.970 112.100 115.970 112.260 ;
        RECT 116.860 112.100 117.860 112.260 ;
        RECT 55.895 111.090 56.895 112.090 ;
        RECT 71.690 111.710 71.940 112.100 ;
        RECT 94.350 111.710 94.600 112.100 ;
        RECT 117.010 111.710 117.260 112.100 ;
        RECT 71.655 111.450 71.975 111.710 ;
        RECT 94.315 111.450 94.635 111.710 ;
        RECT 116.975 111.450 117.295 111.710 ;
        RECT 56.270 109.470 56.520 111.090 ;
        RECT 56.220 107.250 56.570 109.470 ;
        RECT 53.230 104.530 54.230 105.530 ;
        RECT 75.890 104.530 76.890 105.530 ;
        RECT 98.550 104.530 99.550 105.530 ;
        RECT 121.210 104.530 122.210 105.530 ;
        RECT 53.930 104.210 54.180 104.530 ;
        RECT 76.590 104.210 76.840 104.530 ;
        RECT 99.250 104.210 99.500 104.530 ;
        RECT 121.910 104.210 122.160 104.530 ;
        RECT 38.590 101.930 39.590 102.640 ;
        RECT 53.880 101.990 54.230 104.210 ;
        RECT 38.590 101.690 40.060 101.930 ;
        RECT 38.590 101.640 39.590 101.690 ;
        RECT 39.820 95.160 40.060 101.690 ;
        RECT 44.930 95.160 45.930 95.770 ;
        RECT 46.990 95.160 47.990 95.760 ;
        RECT 48.880 95.160 49.880 95.760 ;
        RECT 53.940 95.160 54.180 101.990 ;
        RECT 61.250 101.930 62.250 102.640 ;
        RECT 76.540 101.990 76.890 104.210 ;
        RECT 61.250 101.690 62.720 101.930 ;
        RECT 61.250 101.640 62.250 101.690 ;
        RECT 39.820 94.920 54.180 95.160 ;
        RECT 62.480 95.160 62.720 101.690 ;
        RECT 67.590 95.160 68.590 95.770 ;
        RECT 69.650 95.160 70.650 95.760 ;
        RECT 71.540 95.160 72.540 95.760 ;
        RECT 76.600 95.160 76.840 101.990 ;
        RECT 83.910 101.930 84.910 102.640 ;
        RECT 99.200 101.990 99.550 104.210 ;
        RECT 83.910 101.690 85.380 101.930 ;
        RECT 83.910 101.640 84.910 101.690 ;
        RECT 62.480 94.920 76.840 95.160 ;
        RECT 85.140 95.160 85.380 101.690 ;
        RECT 90.250 95.160 91.250 95.770 ;
        RECT 92.310 95.160 93.310 95.760 ;
        RECT 94.200 95.160 95.200 95.760 ;
        RECT 99.260 95.160 99.500 101.990 ;
        RECT 106.570 101.930 107.570 102.640 ;
        RECT 121.860 101.990 122.210 104.210 ;
        RECT 106.570 101.690 108.040 101.930 ;
        RECT 106.570 101.640 107.570 101.690 ;
        RECT 85.140 94.920 99.500 95.160 ;
        RECT 107.800 95.160 108.040 101.690 ;
        RECT 112.910 95.160 113.910 95.770 ;
        RECT 114.970 95.160 115.970 95.760 ;
        RECT 116.860 95.160 117.860 95.760 ;
        RECT 121.920 95.160 122.160 101.990 ;
        RECT 107.800 94.920 122.160 95.160 ;
        RECT 44.930 94.770 45.930 94.920 ;
        RECT 46.990 94.760 47.990 94.920 ;
        RECT 48.880 94.760 49.880 94.920 ;
        RECT 67.590 94.770 68.590 94.920 ;
        RECT 69.650 94.760 70.650 94.920 ;
        RECT 71.540 94.760 72.540 94.920 ;
        RECT 90.250 94.770 91.250 94.920 ;
        RECT 92.310 94.760 93.310 94.920 ;
        RECT 94.200 94.760 95.200 94.920 ;
        RECT 112.910 94.770 113.910 94.920 ;
        RECT 114.970 94.760 115.970 94.920 ;
        RECT 116.860 94.760 117.860 94.920 ;
        RECT 49.030 94.370 49.280 94.760 ;
        RECT 71.690 94.370 71.940 94.760 ;
        RECT 94.350 94.370 94.600 94.760 ;
        RECT 117.010 94.370 117.260 94.760 ;
        RECT 48.995 94.110 49.315 94.370 ;
        RECT 71.655 94.110 71.975 94.370 ;
        RECT 94.315 94.110 94.635 94.370 ;
        RECT 116.975 94.110 117.295 94.370 ;
        RECT 53.230 87.190 54.230 88.190 ;
        RECT 75.890 87.190 76.890 88.190 ;
        RECT 98.550 87.190 99.550 88.190 ;
        RECT 121.210 87.190 122.210 88.190 ;
        RECT 53.930 86.870 54.180 87.190 ;
        RECT 76.590 86.870 76.840 87.190 ;
        RECT 99.250 86.870 99.500 87.190 ;
        RECT 121.910 86.870 122.160 87.190 ;
        RECT 38.590 84.590 39.590 85.300 ;
        RECT 53.880 84.650 54.230 86.870 ;
        RECT 38.590 84.350 40.060 84.590 ;
        RECT 38.590 84.300 39.590 84.350 ;
        RECT 39.820 77.820 40.060 84.350 ;
        RECT 44.930 77.820 45.930 78.430 ;
        RECT 46.990 77.820 47.990 78.420 ;
        RECT 48.880 77.820 49.880 78.420 ;
        RECT 53.940 77.820 54.180 84.650 ;
        RECT 61.250 84.590 62.250 85.300 ;
        RECT 76.540 84.650 76.890 86.870 ;
        RECT 61.250 84.350 62.720 84.590 ;
        RECT 61.250 84.300 62.250 84.350 ;
        RECT 39.820 77.580 54.180 77.820 ;
        RECT 62.480 77.820 62.720 84.350 ;
        RECT 67.590 77.820 68.590 78.430 ;
        RECT 69.650 77.820 70.650 78.420 ;
        RECT 71.540 77.820 72.540 78.420 ;
        RECT 76.600 77.820 76.840 84.650 ;
        RECT 83.910 84.590 84.910 85.300 ;
        RECT 99.200 84.650 99.550 86.870 ;
        RECT 83.910 84.350 85.380 84.590 ;
        RECT 83.910 84.300 84.910 84.350 ;
        RECT 62.480 77.580 76.840 77.820 ;
        RECT 85.140 77.820 85.380 84.350 ;
        RECT 90.250 77.820 91.250 78.430 ;
        RECT 92.310 77.820 93.310 78.420 ;
        RECT 94.200 77.820 95.200 78.420 ;
        RECT 99.260 77.820 99.500 84.650 ;
        RECT 106.570 84.590 107.570 85.300 ;
        RECT 121.860 84.650 122.210 86.870 ;
        RECT 106.570 84.350 108.040 84.590 ;
        RECT 106.570 84.300 107.570 84.350 ;
        RECT 85.140 77.580 99.500 77.820 ;
        RECT 107.800 77.820 108.040 84.350 ;
        RECT 112.910 77.820 113.910 78.430 ;
        RECT 114.970 77.820 115.970 78.420 ;
        RECT 116.860 77.820 117.860 78.420 ;
        RECT 121.920 77.820 122.160 84.650 ;
        RECT 107.800 77.580 122.160 77.820 ;
        RECT 44.930 77.430 45.930 77.580 ;
        RECT 46.990 77.420 47.990 77.580 ;
        RECT 48.880 77.420 49.880 77.580 ;
        RECT 67.590 77.430 68.590 77.580 ;
        RECT 69.650 77.420 70.650 77.580 ;
        RECT 71.540 77.420 72.540 77.580 ;
        RECT 90.250 77.430 91.250 77.580 ;
        RECT 92.310 77.420 93.310 77.580 ;
        RECT 94.200 77.420 95.200 77.580 ;
        RECT 112.910 77.430 113.910 77.580 ;
        RECT 114.970 77.420 115.970 77.580 ;
        RECT 116.860 77.420 117.860 77.580 ;
        RECT 49.030 77.030 49.280 77.420 ;
        RECT 71.690 77.030 71.940 77.420 ;
        RECT 94.350 77.030 94.600 77.420 ;
        RECT 117.010 77.030 117.260 77.420 ;
        RECT 48.995 76.770 49.315 77.030 ;
        RECT 71.655 76.770 71.975 77.030 ;
        RECT 94.315 76.770 94.635 77.030 ;
        RECT 116.975 76.770 117.295 77.030 ;
        RECT 53.230 69.850 54.230 70.850 ;
        RECT 75.890 69.850 76.890 70.850 ;
        RECT 98.550 69.850 99.550 70.850 ;
        RECT 121.210 69.850 122.210 70.850 ;
        RECT 53.930 69.530 54.180 69.850 ;
        RECT 76.590 69.530 76.840 69.850 ;
        RECT 99.250 69.530 99.500 69.850 ;
        RECT 121.910 69.530 122.160 69.850 ;
        RECT 38.590 67.250 39.590 67.960 ;
        RECT 53.880 67.310 54.230 69.530 ;
        RECT 38.590 67.010 40.060 67.250 ;
        RECT 38.590 66.960 39.590 67.010 ;
        RECT 39.820 60.480 40.060 67.010 ;
        RECT 44.930 60.480 45.930 61.090 ;
        RECT 46.990 60.480 47.990 61.080 ;
        RECT 48.880 60.480 49.880 61.080 ;
        RECT 53.940 60.480 54.180 67.310 ;
        RECT 61.250 67.250 62.250 67.960 ;
        RECT 76.540 67.310 76.890 69.530 ;
        RECT 61.250 67.010 62.720 67.250 ;
        RECT 61.250 66.960 62.250 67.010 ;
        RECT 39.820 60.240 54.180 60.480 ;
        RECT 62.480 60.480 62.720 67.010 ;
        RECT 67.590 60.480 68.590 61.090 ;
        RECT 69.650 60.480 70.650 61.080 ;
        RECT 71.540 60.480 72.540 61.080 ;
        RECT 76.600 60.480 76.840 67.310 ;
        RECT 83.910 67.250 84.910 67.960 ;
        RECT 99.200 67.310 99.550 69.530 ;
        RECT 83.910 67.010 85.380 67.250 ;
        RECT 83.910 66.960 84.910 67.010 ;
        RECT 62.480 60.240 76.840 60.480 ;
        RECT 85.140 60.480 85.380 67.010 ;
        RECT 90.250 60.480 91.250 61.090 ;
        RECT 92.310 60.480 93.310 61.080 ;
        RECT 94.200 60.480 95.200 61.080 ;
        RECT 99.260 60.480 99.500 67.310 ;
        RECT 106.570 67.250 107.570 67.960 ;
        RECT 121.860 67.310 122.210 69.530 ;
        RECT 106.570 67.010 108.040 67.250 ;
        RECT 106.570 66.960 107.570 67.010 ;
        RECT 85.140 60.240 99.500 60.480 ;
        RECT 107.800 60.480 108.040 67.010 ;
        RECT 112.910 60.480 113.910 61.090 ;
        RECT 114.970 60.480 115.970 61.080 ;
        RECT 116.860 60.480 117.860 61.080 ;
        RECT 121.920 60.480 122.160 67.310 ;
        RECT 107.800 60.240 122.160 60.480 ;
        RECT 44.930 60.090 45.930 60.240 ;
        RECT 46.990 60.080 47.990 60.240 ;
        RECT 48.880 60.080 49.880 60.240 ;
        RECT 67.590 60.090 68.590 60.240 ;
        RECT 69.650 60.080 70.650 60.240 ;
        RECT 71.540 60.080 72.540 60.240 ;
        RECT 90.250 60.090 91.250 60.240 ;
        RECT 92.310 60.080 93.310 60.240 ;
        RECT 94.200 60.080 95.200 60.240 ;
        RECT 112.910 60.090 113.910 60.240 ;
        RECT 114.970 60.080 115.970 60.240 ;
        RECT 116.860 60.080 117.860 60.240 ;
        RECT 49.030 59.690 49.280 60.080 ;
        RECT 71.690 59.690 71.940 60.080 ;
        RECT 94.350 59.690 94.600 60.080 ;
        RECT 117.010 59.690 117.260 60.080 ;
        RECT 48.995 59.430 49.315 59.690 ;
        RECT 71.655 59.430 71.975 59.690 ;
        RECT 94.315 59.430 94.635 59.690 ;
        RECT 116.975 59.430 117.295 59.690 ;
        RECT 53.230 51.850 54.230 52.850 ;
        RECT 75.890 51.850 76.890 52.850 ;
        RECT 98.550 51.850 99.550 52.850 ;
        RECT 121.210 51.850 122.210 52.850 ;
        RECT 53.930 51.530 54.180 51.850 ;
        RECT 76.590 51.530 76.840 51.850 ;
        RECT 99.250 51.530 99.500 51.850 ;
        RECT 121.910 51.530 122.160 51.850 ;
        RECT 53.880 49.310 54.230 51.530 ;
        RECT 76.540 49.310 76.890 51.530 ;
        RECT 99.200 49.310 99.550 51.530 ;
        RECT 121.860 49.310 122.210 51.530 ;
        RECT 44.930 42.480 45.930 43.090 ;
        RECT 46.990 42.480 47.990 43.080 ;
        RECT 48.880 42.480 49.880 43.080 ;
        RECT 53.940 42.480 54.180 49.310 ;
        RECT 44.930 42.240 54.180 42.480 ;
        RECT 67.590 42.480 68.590 43.090 ;
        RECT 69.650 42.480 70.650 43.080 ;
        RECT 71.540 42.480 72.540 43.080 ;
        RECT 76.600 42.480 76.840 49.310 ;
        RECT 67.590 42.240 76.840 42.480 ;
        RECT 90.250 42.480 91.250 43.090 ;
        RECT 92.310 42.480 93.310 43.080 ;
        RECT 94.200 42.480 95.200 43.080 ;
        RECT 99.260 42.480 99.500 49.310 ;
        RECT 90.250 42.240 99.500 42.480 ;
        RECT 112.910 42.480 113.910 43.090 ;
        RECT 114.970 42.480 115.970 43.080 ;
        RECT 116.860 42.480 117.860 43.080 ;
        RECT 121.920 42.480 122.160 49.310 ;
        RECT 125.830 46.125 126.830 116.215 ;
        RECT 112.910 42.240 122.160 42.480 ;
        RECT 44.930 42.090 45.930 42.240 ;
        RECT 46.990 42.080 47.990 42.240 ;
        RECT 48.880 42.080 49.880 42.240 ;
        RECT 67.590 42.090 68.590 42.240 ;
        RECT 69.650 42.080 70.650 42.240 ;
        RECT 71.540 42.080 72.540 42.240 ;
        RECT 90.250 42.090 91.250 42.240 ;
        RECT 92.310 42.080 93.310 42.240 ;
        RECT 94.200 42.080 95.200 42.240 ;
        RECT 112.910 42.090 113.910 42.240 ;
        RECT 114.970 42.080 115.970 42.240 ;
        RECT 116.860 42.080 117.860 42.240 ;
        RECT 49.030 41.690 49.280 42.080 ;
        RECT 71.690 41.690 71.940 42.080 ;
        RECT 94.350 41.690 94.600 42.080 ;
        RECT 117.010 41.690 117.260 42.080 ;
        RECT 48.995 41.430 49.315 41.690 ;
        RECT 71.655 41.430 71.975 41.690 ;
        RECT 94.315 41.430 94.635 41.690 ;
        RECT 116.975 41.430 117.295 41.690 ;
      LAYER via2 ;
        RECT 50.295 186.450 50.575 186.730 ;
        RECT 50.695 186.450 50.975 186.730 ;
        RECT 51.095 186.450 51.375 186.730 ;
        RECT 51.495 186.450 51.775 186.730 ;
        RECT 68.805 186.450 69.085 186.730 ;
        RECT 69.205 186.450 69.485 186.730 ;
        RECT 69.605 186.450 69.885 186.730 ;
        RECT 70.005 186.450 70.285 186.730 ;
        RECT 87.315 186.450 87.595 186.730 ;
        RECT 87.715 186.450 87.995 186.730 ;
        RECT 88.115 186.450 88.395 186.730 ;
        RECT 88.515 186.450 88.795 186.730 ;
        RECT 105.825 186.450 106.105 186.730 ;
        RECT 106.225 186.450 106.505 186.730 ;
        RECT 106.625 186.450 106.905 186.730 ;
        RECT 107.025 186.450 107.305 186.730 ;
        RECT 50.295 181.010 50.575 181.290 ;
        RECT 50.695 181.010 50.975 181.290 ;
        RECT 51.095 181.010 51.375 181.290 ;
        RECT 51.495 181.010 51.775 181.290 ;
        RECT 68.805 181.010 69.085 181.290 ;
        RECT 69.205 181.010 69.485 181.290 ;
        RECT 69.605 181.010 69.885 181.290 ;
        RECT 70.005 181.010 70.285 181.290 ;
        RECT 87.315 181.010 87.595 181.290 ;
        RECT 87.715 181.010 87.995 181.290 ;
        RECT 88.115 181.010 88.395 181.290 ;
        RECT 88.515 181.010 88.795 181.290 ;
        RECT 105.825 181.010 106.105 181.290 ;
        RECT 106.225 181.010 106.505 181.290 ;
        RECT 106.625 181.010 106.905 181.290 ;
        RECT 107.025 181.010 107.305 181.290 ;
        RECT 50.295 175.570 50.575 175.850 ;
        RECT 50.695 175.570 50.975 175.850 ;
        RECT 51.095 175.570 51.375 175.850 ;
        RECT 51.495 175.570 51.775 175.850 ;
        RECT 68.805 175.570 69.085 175.850 ;
        RECT 69.205 175.570 69.485 175.850 ;
        RECT 69.605 175.570 69.885 175.850 ;
        RECT 70.005 175.570 70.285 175.850 ;
        RECT 87.315 175.570 87.595 175.850 ;
        RECT 87.715 175.570 87.995 175.850 ;
        RECT 88.115 175.570 88.395 175.850 ;
        RECT 88.515 175.570 88.795 175.850 ;
        RECT 105.825 175.570 106.105 175.850 ;
        RECT 106.225 175.570 106.505 175.850 ;
        RECT 106.625 175.570 106.905 175.850 ;
        RECT 107.025 175.570 107.305 175.850 ;
        RECT 50.295 170.130 50.575 170.410 ;
        RECT 50.695 170.130 50.975 170.410 ;
        RECT 51.095 170.130 51.375 170.410 ;
        RECT 51.495 170.130 51.775 170.410 ;
        RECT 68.805 170.130 69.085 170.410 ;
        RECT 69.205 170.130 69.485 170.410 ;
        RECT 69.605 170.130 69.885 170.410 ;
        RECT 70.005 170.130 70.285 170.410 ;
        RECT 87.315 170.130 87.595 170.410 ;
        RECT 87.715 170.130 87.995 170.410 ;
        RECT 88.115 170.130 88.395 170.410 ;
        RECT 88.515 170.130 88.795 170.410 ;
        RECT 105.825 170.130 106.105 170.410 ;
        RECT 106.225 170.130 106.505 170.410 ;
        RECT 106.625 170.130 106.905 170.410 ;
        RECT 107.025 170.130 107.305 170.410 ;
        RECT 50.295 164.690 50.575 164.970 ;
        RECT 50.695 164.690 50.975 164.970 ;
        RECT 51.095 164.690 51.375 164.970 ;
        RECT 51.495 164.690 51.775 164.970 ;
        RECT 68.805 164.690 69.085 164.970 ;
        RECT 69.205 164.690 69.485 164.970 ;
        RECT 69.605 164.690 69.885 164.970 ;
        RECT 70.005 164.690 70.285 164.970 ;
        RECT 87.315 164.690 87.595 164.970 ;
        RECT 87.715 164.690 87.995 164.970 ;
        RECT 88.115 164.690 88.395 164.970 ;
        RECT 88.515 164.690 88.795 164.970 ;
        RECT 105.825 164.690 106.105 164.970 ;
        RECT 106.225 164.690 106.505 164.970 ;
        RECT 106.625 164.690 106.905 164.970 ;
        RECT 107.025 164.690 107.305 164.970 ;
        RECT 50.295 159.250 50.575 159.530 ;
        RECT 50.695 159.250 50.975 159.530 ;
        RECT 51.095 159.250 51.375 159.530 ;
        RECT 51.495 159.250 51.775 159.530 ;
        RECT 68.805 159.250 69.085 159.530 ;
        RECT 69.205 159.250 69.485 159.530 ;
        RECT 69.605 159.250 69.885 159.530 ;
        RECT 70.005 159.250 70.285 159.530 ;
        RECT 87.315 159.250 87.595 159.530 ;
        RECT 87.715 159.250 87.995 159.530 ;
        RECT 88.115 159.250 88.395 159.530 ;
        RECT 88.515 159.250 88.795 159.530 ;
        RECT 105.825 159.250 106.105 159.530 ;
        RECT 106.225 159.250 106.505 159.530 ;
        RECT 106.625 159.250 106.905 159.530 ;
        RECT 107.025 159.250 107.305 159.530 ;
        RECT 75.940 121.920 76.840 122.820 ;
        RECT 98.600 121.920 99.500 122.820 ;
        RECT 121.260 121.920 122.160 122.820 ;
        RECT 61.300 119.030 62.200 119.930 ;
        RECT 32.920 116.200 33.920 117.200 ;
        RECT 67.640 112.160 68.540 113.060 ;
        RECT 69.700 112.150 70.600 113.050 ;
        RECT 71.590 112.150 72.490 113.050 ;
        RECT 83.960 119.030 84.860 119.930 ;
        RECT 90.300 112.160 91.200 113.060 ;
        RECT 92.360 112.150 93.260 113.050 ;
        RECT 94.250 112.150 95.150 113.050 ;
        RECT 106.620 119.030 107.520 119.930 ;
        RECT 112.960 112.160 113.860 113.060 ;
        RECT 115.020 112.150 115.920 113.050 ;
        RECT 116.910 112.150 117.810 113.050 ;
        RECT 125.855 116.215 126.805 117.165 ;
        RECT 55.945 111.140 56.845 112.040 ;
        RECT 53.280 104.580 54.180 105.480 ;
        RECT 75.940 104.580 76.840 105.480 ;
        RECT 98.600 104.580 99.500 105.480 ;
        RECT 121.260 104.580 122.160 105.480 ;
        RECT 38.640 101.690 39.540 102.590 ;
        RECT 32.920 98.850 33.920 99.850 ;
        RECT 44.980 94.820 45.880 95.720 ;
        RECT 47.040 94.810 47.940 95.710 ;
        RECT 48.930 94.810 49.830 95.710 ;
        RECT 61.300 101.690 62.200 102.590 ;
        RECT 67.640 94.820 68.540 95.720 ;
        RECT 69.700 94.810 70.600 95.710 ;
        RECT 71.590 94.810 72.490 95.710 ;
        RECT 83.960 101.690 84.860 102.590 ;
        RECT 90.300 94.820 91.200 95.720 ;
        RECT 92.360 94.810 93.260 95.710 ;
        RECT 94.250 94.810 95.150 95.710 ;
        RECT 106.620 101.690 107.520 102.590 ;
        RECT 112.960 94.820 113.860 95.720 ;
        RECT 115.020 94.810 115.920 95.710 ;
        RECT 116.910 94.810 117.810 95.710 ;
        RECT 125.830 98.850 126.830 99.850 ;
        RECT 53.280 87.240 54.180 88.140 ;
        RECT 75.940 87.240 76.840 88.140 ;
        RECT 98.600 87.240 99.500 88.140 ;
        RECT 121.260 87.240 122.160 88.140 ;
        RECT 38.640 84.350 39.540 85.250 ;
        RECT 32.920 81.510 33.920 82.510 ;
        RECT 44.980 77.480 45.880 78.380 ;
        RECT 47.040 77.470 47.940 78.370 ;
        RECT 48.930 77.470 49.830 78.370 ;
        RECT 61.300 84.350 62.200 85.250 ;
        RECT 67.640 77.480 68.540 78.380 ;
        RECT 69.700 77.470 70.600 78.370 ;
        RECT 71.590 77.470 72.490 78.370 ;
        RECT 83.960 84.350 84.860 85.250 ;
        RECT 90.300 77.480 91.200 78.380 ;
        RECT 92.360 77.470 93.260 78.370 ;
        RECT 94.250 77.470 95.150 78.370 ;
        RECT 106.620 84.350 107.520 85.250 ;
        RECT 112.960 77.480 113.860 78.380 ;
        RECT 115.020 77.470 115.920 78.370 ;
        RECT 116.910 77.470 117.810 78.370 ;
        RECT 125.830 81.500 126.830 82.500 ;
        RECT 53.280 69.900 54.180 70.800 ;
        RECT 75.940 69.900 76.840 70.800 ;
        RECT 98.600 69.900 99.500 70.800 ;
        RECT 121.260 69.900 122.160 70.800 ;
        RECT 38.640 67.010 39.540 67.910 ;
        RECT 32.945 64.195 33.895 65.145 ;
        RECT 44.980 60.140 45.880 61.040 ;
        RECT 47.040 60.130 47.940 61.030 ;
        RECT 48.930 60.130 49.830 61.030 ;
        RECT 61.300 67.010 62.200 67.910 ;
        RECT 67.640 60.140 68.540 61.040 ;
        RECT 69.700 60.130 70.600 61.030 ;
        RECT 71.590 60.130 72.490 61.030 ;
        RECT 83.960 67.010 84.860 67.910 ;
        RECT 90.300 60.140 91.200 61.040 ;
        RECT 92.360 60.130 93.260 61.030 ;
        RECT 94.250 60.130 95.150 61.030 ;
        RECT 106.620 67.010 107.520 67.910 ;
        RECT 112.960 60.140 113.860 61.040 ;
        RECT 115.020 60.130 115.920 61.030 ;
        RECT 116.910 60.130 117.810 61.030 ;
        RECT 125.830 64.170 126.830 65.170 ;
        RECT 53.280 51.900 54.180 52.800 ;
        RECT 75.940 51.900 76.840 52.800 ;
        RECT 98.600 51.900 99.500 52.800 ;
        RECT 121.260 51.900 122.160 52.800 ;
        RECT 32.920 46.170 33.920 47.170 ;
        RECT 44.980 42.140 45.880 43.040 ;
        RECT 47.040 42.130 47.940 43.030 ;
        RECT 48.930 42.130 49.830 43.030 ;
        RECT 67.640 42.140 68.540 43.040 ;
        RECT 69.700 42.130 70.600 43.030 ;
        RECT 71.590 42.130 72.490 43.030 ;
        RECT 90.300 42.140 91.200 43.040 ;
        RECT 92.360 42.130 93.260 43.030 ;
        RECT 94.250 42.130 95.150 43.030 ;
        RECT 112.960 42.140 113.860 43.040 ;
        RECT 115.020 42.130 115.920 43.030 ;
        RECT 116.910 42.130 117.810 43.030 ;
        RECT 125.830 46.170 126.830 47.170 ;
      LAYER met3 ;
        RECT 50.245 186.425 51.825 186.755 ;
        RECT 68.755 186.425 70.335 186.755 ;
        RECT 87.265 186.425 88.845 186.755 ;
        RECT 105.775 186.425 107.355 186.755 ;
        RECT 50.245 180.985 51.825 181.315 ;
        RECT 68.755 180.985 70.335 181.315 ;
        RECT 87.265 180.985 88.845 181.315 ;
        RECT 105.775 180.985 107.355 181.315 ;
        RECT 50.245 175.545 51.825 175.875 ;
        RECT 68.755 175.545 70.335 175.875 ;
        RECT 87.265 175.545 88.845 175.875 ;
        RECT 105.775 175.545 107.355 175.875 ;
        RECT 50.245 170.105 51.825 170.435 ;
        RECT 68.755 170.105 70.335 170.435 ;
        RECT 87.265 170.105 88.845 170.435 ;
        RECT 105.775 170.105 107.355 170.435 ;
        RECT 50.245 164.665 51.825 164.995 ;
        RECT 68.755 164.665 70.335 164.995 ;
        RECT 87.265 164.665 88.845 164.995 ;
        RECT 105.775 164.665 107.355 164.995 ;
        RECT 50.245 159.225 51.825 159.555 ;
        RECT 68.755 159.225 70.335 159.555 ;
        RECT 87.265 159.225 88.845 159.555 ;
        RECT 105.775 159.225 107.355 159.555 ;
        RECT 12.000 137.000 116.620 138.600 ;
        RECT 32.895 117.190 33.945 117.225 ;
        RECT 61.250 117.190 62.250 119.980 ;
        RECT 75.890 117.190 76.890 122.870 ;
        RECT 83.910 117.190 84.910 119.980 ;
        RECT 98.550 117.190 99.550 122.870 ;
        RECT 106.570 117.190 107.570 119.980 ;
        RECT 121.210 117.190 122.210 122.870 ;
        RECT 30.890 117.180 128.830 117.190 ;
        RECT 30.880 116.180 128.840 117.180 ;
        RECT 32.895 116.175 33.945 116.180 ;
        RECT 55.895 111.090 56.895 116.180 ;
        RECT 67.590 112.110 68.590 116.180 ;
        RECT 69.650 112.100 70.650 116.180 ;
        RECT 71.540 112.100 72.540 116.180 ;
        RECT 90.250 112.110 91.250 116.180 ;
        RECT 92.310 112.100 93.310 116.180 ;
        RECT 94.200 112.100 95.200 116.180 ;
        RECT 112.910 112.110 113.910 116.180 ;
        RECT 114.970 112.100 115.970 116.180 ;
        RECT 116.860 112.100 117.860 116.180 ;
        RECT 32.895 99.850 33.945 99.875 ;
        RECT 38.590 99.850 39.590 102.640 ;
        RECT 53.230 99.850 54.230 105.530 ;
        RECT 61.250 99.850 62.250 102.640 ;
        RECT 75.890 99.850 76.890 105.530 ;
        RECT 83.910 99.850 84.910 102.640 ;
        RECT 98.550 99.850 99.550 105.530 ;
        RECT 106.570 99.850 107.570 102.640 ;
        RECT 121.210 99.850 122.210 105.530 ;
        RECT 125.805 99.850 126.855 99.875 ;
        RECT 30.890 99.840 128.830 99.850 ;
        RECT 30.880 98.840 128.840 99.840 ;
        RECT 32.895 98.825 33.945 98.840 ;
        RECT 44.930 94.770 45.930 98.840 ;
        RECT 46.990 94.760 47.990 98.840 ;
        RECT 48.880 94.760 49.880 98.840 ;
        RECT 67.590 94.770 68.590 98.840 ;
        RECT 69.650 94.760 70.650 98.840 ;
        RECT 71.540 94.760 72.540 98.840 ;
        RECT 90.250 94.770 91.250 98.840 ;
        RECT 92.310 94.760 93.310 98.840 ;
        RECT 94.200 94.760 95.200 98.840 ;
        RECT 112.910 94.770 113.910 98.840 ;
        RECT 114.970 94.760 115.970 98.840 ;
        RECT 116.860 94.760 117.860 98.840 ;
        RECT 125.805 98.825 126.855 98.840 ;
        RECT 32.895 82.510 33.945 82.535 ;
        RECT 38.590 82.510 39.590 85.300 ;
        RECT 53.230 82.510 54.230 88.190 ;
        RECT 61.250 82.510 62.250 85.300 ;
        RECT 75.890 82.510 76.890 88.190 ;
        RECT 83.910 82.510 84.910 85.300 ;
        RECT 98.550 82.510 99.550 88.190 ;
        RECT 106.570 82.510 107.570 85.300 ;
        RECT 121.210 82.510 122.210 88.190 ;
        RECT 125.805 82.510 126.855 82.525 ;
        RECT 30.890 82.500 128.830 82.510 ;
        RECT 30.880 81.500 128.840 82.500 ;
        RECT 32.895 81.485 33.945 81.500 ;
        RECT 44.930 77.430 45.930 81.500 ;
        RECT 46.990 77.420 47.990 81.500 ;
        RECT 48.880 77.420 49.880 81.500 ;
        RECT 67.590 77.430 68.590 81.500 ;
        RECT 69.650 77.420 70.650 81.500 ;
        RECT 71.540 77.420 72.540 81.500 ;
        RECT 90.250 77.430 91.250 81.500 ;
        RECT 92.310 77.420 93.310 81.500 ;
        RECT 94.200 77.420 95.200 81.500 ;
        RECT 112.910 77.430 113.910 81.500 ;
        RECT 114.970 77.420 115.970 81.500 ;
        RECT 116.860 77.420 117.860 81.500 ;
        RECT 125.805 81.475 126.855 81.500 ;
        RECT 38.590 65.170 39.590 67.960 ;
        RECT 53.230 65.170 54.230 70.850 ;
        RECT 61.250 65.170 62.250 67.960 ;
        RECT 75.890 65.170 76.890 70.850 ;
        RECT 83.910 65.170 84.910 67.960 ;
        RECT 98.550 65.170 99.550 70.850 ;
        RECT 106.570 65.170 107.570 67.960 ;
        RECT 121.210 65.170 122.210 70.850 ;
        RECT 125.805 65.170 126.855 65.195 ;
        RECT 30.890 65.160 128.830 65.170 ;
        RECT 30.880 64.160 128.840 65.160 ;
        RECT 44.930 60.090 45.930 64.160 ;
        RECT 46.990 60.080 47.990 64.160 ;
        RECT 48.880 60.080 49.880 64.160 ;
        RECT 67.590 60.090 68.590 64.160 ;
        RECT 69.650 60.080 70.650 64.160 ;
        RECT 71.540 60.080 72.540 64.160 ;
        RECT 90.250 60.090 91.250 64.160 ;
        RECT 92.310 60.080 93.310 64.160 ;
        RECT 94.200 60.080 95.200 64.160 ;
        RECT 112.910 60.090 113.910 64.160 ;
        RECT 114.970 60.080 115.970 64.160 ;
        RECT 116.860 60.080 117.860 64.160 ;
        RECT 125.805 64.145 126.855 64.160 ;
        RECT 32.895 47.170 33.945 47.195 ;
        RECT 53.230 47.170 54.230 52.850 ;
        RECT 75.890 47.170 76.890 52.850 ;
        RECT 98.550 47.170 99.550 52.850 ;
        RECT 121.210 47.170 122.210 52.850 ;
        RECT 125.805 47.170 126.855 47.195 ;
        RECT 30.890 47.160 128.830 47.170 ;
        RECT 30.880 46.160 128.840 47.160 ;
        RECT 32.895 46.145 33.945 46.160 ;
        RECT 44.930 42.090 45.930 46.160 ;
        RECT 46.990 42.080 47.990 46.160 ;
        RECT 48.880 42.080 49.880 46.160 ;
        RECT 67.590 42.090 68.590 46.160 ;
        RECT 69.650 42.080 70.650 46.160 ;
        RECT 71.540 42.080 72.540 46.160 ;
        RECT 90.250 42.090 91.250 46.160 ;
        RECT 92.310 42.080 93.310 46.160 ;
        RECT 94.200 42.080 95.200 46.160 ;
        RECT 112.910 42.090 113.910 46.160 ;
        RECT 114.970 42.080 115.970 46.160 ;
        RECT 116.860 42.080 117.860 46.160 ;
        RECT 125.805 46.145 126.855 46.160 ;
      LAYER via3 ;
        RECT 50.275 186.430 50.595 186.750 ;
        RECT 50.675 186.430 50.995 186.750 ;
        RECT 51.075 186.430 51.395 186.750 ;
        RECT 51.475 186.430 51.795 186.750 ;
        RECT 68.785 186.430 69.105 186.750 ;
        RECT 69.185 186.430 69.505 186.750 ;
        RECT 69.585 186.430 69.905 186.750 ;
        RECT 69.985 186.430 70.305 186.750 ;
        RECT 87.295 186.430 87.615 186.750 ;
        RECT 87.695 186.430 88.015 186.750 ;
        RECT 88.095 186.430 88.415 186.750 ;
        RECT 88.495 186.430 88.815 186.750 ;
        RECT 105.805 186.430 106.125 186.750 ;
        RECT 106.205 186.430 106.525 186.750 ;
        RECT 106.605 186.430 106.925 186.750 ;
        RECT 107.005 186.430 107.325 186.750 ;
        RECT 50.275 180.990 50.595 181.310 ;
        RECT 50.675 180.990 50.995 181.310 ;
        RECT 51.075 180.990 51.395 181.310 ;
        RECT 51.475 180.990 51.795 181.310 ;
        RECT 68.785 180.990 69.105 181.310 ;
        RECT 69.185 180.990 69.505 181.310 ;
        RECT 69.585 180.990 69.905 181.310 ;
        RECT 69.985 180.990 70.305 181.310 ;
        RECT 87.295 180.990 87.615 181.310 ;
        RECT 87.695 180.990 88.015 181.310 ;
        RECT 88.095 180.990 88.415 181.310 ;
        RECT 88.495 180.990 88.815 181.310 ;
        RECT 105.805 180.990 106.125 181.310 ;
        RECT 106.205 180.990 106.525 181.310 ;
        RECT 106.605 180.990 106.925 181.310 ;
        RECT 107.005 180.990 107.325 181.310 ;
        RECT 50.275 175.550 50.595 175.870 ;
        RECT 50.675 175.550 50.995 175.870 ;
        RECT 51.075 175.550 51.395 175.870 ;
        RECT 51.475 175.550 51.795 175.870 ;
        RECT 68.785 175.550 69.105 175.870 ;
        RECT 69.185 175.550 69.505 175.870 ;
        RECT 69.585 175.550 69.905 175.870 ;
        RECT 69.985 175.550 70.305 175.870 ;
        RECT 87.295 175.550 87.615 175.870 ;
        RECT 87.695 175.550 88.015 175.870 ;
        RECT 88.095 175.550 88.415 175.870 ;
        RECT 88.495 175.550 88.815 175.870 ;
        RECT 105.805 175.550 106.125 175.870 ;
        RECT 106.205 175.550 106.525 175.870 ;
        RECT 106.605 175.550 106.925 175.870 ;
        RECT 107.005 175.550 107.325 175.870 ;
        RECT 50.275 170.110 50.595 170.430 ;
        RECT 50.675 170.110 50.995 170.430 ;
        RECT 51.075 170.110 51.395 170.430 ;
        RECT 51.475 170.110 51.795 170.430 ;
        RECT 68.785 170.110 69.105 170.430 ;
        RECT 69.185 170.110 69.505 170.430 ;
        RECT 69.585 170.110 69.905 170.430 ;
        RECT 69.985 170.110 70.305 170.430 ;
        RECT 87.295 170.110 87.615 170.430 ;
        RECT 87.695 170.110 88.015 170.430 ;
        RECT 88.095 170.110 88.415 170.430 ;
        RECT 88.495 170.110 88.815 170.430 ;
        RECT 105.805 170.110 106.125 170.430 ;
        RECT 106.205 170.110 106.525 170.430 ;
        RECT 106.605 170.110 106.925 170.430 ;
        RECT 107.005 170.110 107.325 170.430 ;
        RECT 50.275 164.670 50.595 164.990 ;
        RECT 50.675 164.670 50.995 164.990 ;
        RECT 51.075 164.670 51.395 164.990 ;
        RECT 51.475 164.670 51.795 164.990 ;
        RECT 68.785 164.670 69.105 164.990 ;
        RECT 69.185 164.670 69.505 164.990 ;
        RECT 69.585 164.670 69.905 164.990 ;
        RECT 69.985 164.670 70.305 164.990 ;
        RECT 87.295 164.670 87.615 164.990 ;
        RECT 87.695 164.670 88.015 164.990 ;
        RECT 88.095 164.670 88.415 164.990 ;
        RECT 88.495 164.670 88.815 164.990 ;
        RECT 105.805 164.670 106.125 164.990 ;
        RECT 106.205 164.670 106.525 164.990 ;
        RECT 106.605 164.670 106.925 164.990 ;
        RECT 107.005 164.670 107.325 164.990 ;
        RECT 50.275 159.230 50.595 159.550 ;
        RECT 50.675 159.230 50.995 159.550 ;
        RECT 51.075 159.230 51.395 159.550 ;
        RECT 51.475 159.230 51.795 159.550 ;
        RECT 68.785 159.230 69.105 159.550 ;
        RECT 69.185 159.230 69.505 159.550 ;
        RECT 69.585 159.230 69.905 159.550 ;
        RECT 69.985 159.230 70.305 159.550 ;
        RECT 87.295 159.230 87.615 159.550 ;
        RECT 87.695 159.230 88.015 159.550 ;
        RECT 88.095 159.230 88.415 159.550 ;
        RECT 88.495 159.230 88.815 159.550 ;
        RECT 105.805 159.230 106.125 159.550 ;
        RECT 106.205 159.230 106.525 159.550 ;
        RECT 106.605 159.230 106.925 159.550 ;
        RECT 107.005 159.230 107.325 159.550 ;
        RECT 12.100 137.100 13.500 138.500 ;
        RECT 50.335 137.100 51.735 138.500 ;
        RECT 68.855 137.100 70.255 138.500 ;
        RECT 87.365 137.100 88.765 138.500 ;
        RECT 105.875 137.100 107.275 138.500 ;
        RECT 50.335 116.280 51.735 117.090 ;
        RECT 68.845 116.280 70.245 117.090 ;
        RECT 87.355 116.280 88.755 117.090 ;
        RECT 105.865 116.280 107.265 117.090 ;
        RECT 50.335 98.940 51.735 99.750 ;
        RECT 68.845 98.940 70.245 99.750 ;
        RECT 87.355 98.940 88.755 99.750 ;
        RECT 105.865 98.940 107.265 99.750 ;
        RECT 50.335 81.600 51.735 82.410 ;
        RECT 68.845 81.600 70.245 82.410 ;
        RECT 87.355 81.600 88.755 82.410 ;
        RECT 105.865 81.600 107.265 82.410 ;
        RECT 50.335 64.260 51.735 65.070 ;
        RECT 68.845 64.260 70.245 65.070 ;
        RECT 87.355 64.260 88.755 65.070 ;
        RECT 105.865 64.260 107.265 65.070 ;
        RECT 50.335 46.260 51.735 47.070 ;
        RECT 68.845 46.260 70.245 47.070 ;
        RECT 87.355 46.260 88.755 47.070 ;
        RECT 105.865 46.260 107.265 47.070 ;
      LAYER met4 ;
        RECT 12.000 5.000 13.600 220.760 ;
        RECT 50.235 44.400 51.835 186.850 ;
        RECT 68.745 44.400 70.345 186.850 ;
        RECT 87.255 44.400 88.855 186.850 ;
        RECT 105.765 44.400 107.365 186.850 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 54.675 184.060 55.105 184.845 ;
        RECT 67.555 184.060 67.985 184.845 ;
        RECT 80.435 184.060 80.865 184.845 ;
        RECT 93.315 184.060 93.745 184.845 ;
        RECT 106.195 184.060 106.625 184.845 ;
        RECT 67.555 182.895 67.985 183.680 ;
        RECT 93.315 182.895 93.745 183.680 ;
        RECT 54.675 178.620 55.105 179.405 ;
        RECT 80.435 178.620 80.865 179.405 ;
        RECT 106.195 178.620 106.625 179.405 ;
        RECT 67.555 177.455 67.985 178.240 ;
        RECT 93.315 177.455 93.745 178.240 ;
        RECT 54.675 173.180 55.105 173.965 ;
        RECT 80.435 173.180 80.865 173.965 ;
        RECT 106.195 173.180 106.625 173.965 ;
        RECT 67.555 172.015 67.985 172.800 ;
        RECT 93.315 172.015 93.745 172.800 ;
        RECT 54.675 167.740 55.105 168.525 ;
        RECT 80.435 167.740 80.865 168.525 ;
        RECT 106.195 167.740 106.625 168.525 ;
        RECT 67.555 166.575 67.985 167.360 ;
        RECT 93.315 166.575 93.745 167.360 ;
        RECT 54.675 162.300 55.105 163.085 ;
        RECT 80.435 162.300 80.865 163.085 ;
        RECT 106.195 162.300 106.625 163.085 ;
        RECT 67.555 161.135 67.985 161.920 ;
        RECT 93.315 161.135 93.745 161.920 ;
        RECT 54.675 156.860 55.105 157.645 ;
        RECT 67.555 156.860 67.985 157.645 ;
        RECT 80.435 156.860 80.865 157.645 ;
        RECT 93.315 156.860 93.745 157.645 ;
        RECT 106.195 156.860 106.625 157.645 ;
      LAYER li1 ;
        RECT 41.865 184.705 42.385 185.245 ;
        RECT 41.865 183.955 43.075 184.705 ;
        RECT 44.635 183.955 44.910 184.435 ;
        RECT 45.555 183.955 45.810 184.435 ;
        RECT 46.415 183.955 46.695 184.435 ;
        RECT 48.320 183.955 48.650 184.335 ;
        RECT 49.250 183.955 49.510 184.795 ;
        RECT 50.620 183.955 50.950 184.335 ;
        RECT 51.550 183.955 51.810 184.795 ;
        RECT 52.460 183.955 52.790 184.335 ;
        RECT 53.390 183.955 53.650 184.795 ;
        RECT 54.745 183.955 55.035 184.680 ;
        RECT 55.210 183.955 55.470 184.795 ;
        RECT 56.070 183.955 56.400 184.335 ;
        RECT 57.980 183.955 58.310 184.335 ;
        RECT 58.910 183.955 59.170 184.795 ;
        RECT 59.820 183.955 60.150 184.335 ;
        RECT 60.750 183.955 61.010 184.795 ;
        RECT 61.190 183.955 61.450 184.795 ;
        RECT 62.050 183.955 62.380 184.335 ;
        RECT 63.495 183.955 63.770 184.435 ;
        RECT 64.415 183.955 64.670 184.435 ;
        RECT 65.275 183.955 65.555 184.435 ;
        RECT 66.260 183.955 66.590 184.335 ;
        RECT 67.190 183.955 67.450 184.795 ;
        RECT 67.625 183.955 67.915 184.680 ;
        RECT 68.090 183.955 68.350 184.795 ;
        RECT 68.950 183.955 69.280 184.335 ;
        RECT 70.400 183.955 70.730 184.335 ;
        RECT 71.330 183.955 71.590 184.795 ;
        RECT 71.770 183.955 72.030 184.795 ;
        RECT 72.630 183.955 72.960 184.335 ;
        RECT 74.530 183.955 74.790 184.795 ;
        RECT 75.390 183.955 75.720 184.335 ;
        RECT 76.830 183.955 77.090 184.795 ;
        RECT 78.665 184.725 79.415 185.245 ;
        RECT 77.690 183.955 78.020 184.335 ;
        RECT 78.665 183.955 80.335 184.725 ;
        RECT 80.505 183.955 80.795 184.680 ;
        RECT 82.035 183.955 82.365 184.755 ;
        RECT 82.875 183.955 83.205 184.435 ;
        RECT 83.795 183.955 84.035 184.435 ;
        RECT 84.705 183.955 84.985 184.435 ;
        RECT 85.590 183.955 85.845 184.435 ;
        RECT 86.490 183.955 86.765 184.435 ;
        RECT 87.845 183.955 88.175 184.335 ;
        RECT 89.685 183.955 90.015 184.335 ;
        RECT 91.525 183.955 91.855 184.335 ;
        RECT 93.385 183.955 93.675 184.680 ;
        RECT 93.855 183.955 94.185 184.755 ;
        RECT 94.695 183.955 95.025 184.435 ;
        RECT 95.535 183.955 95.865 184.435 ;
        RECT 96.455 183.955 96.625 184.435 ;
        RECT 97.295 183.955 97.465 184.435 ;
        RECT 98.965 183.955 99.245 184.435 ;
        RECT 99.850 183.955 100.105 184.435 ;
        RECT 100.750 183.955 101.025 184.435 ;
        RECT 102.405 183.955 102.915 184.490 ;
        RECT 104.875 183.955 105.205 184.355 ;
        RECT 106.265 183.955 106.555 184.680 ;
        RECT 107.650 183.955 107.910 184.795 ;
        RECT 115.235 184.705 115.755 185.245 ;
        RECT 108.510 183.955 108.840 184.335 ;
        RECT 109.915 183.955 110.245 184.355 ;
        RECT 112.205 183.955 112.715 184.490 ;
        RECT 114.545 183.955 115.755 184.705 ;
        RECT 41.780 183.785 115.840 183.955 ;
        RECT 41.865 183.035 43.075 183.785 ;
        RECT 41.865 182.495 42.385 183.035 ;
        RECT 44.170 182.945 44.430 183.785 ;
        RECT 45.030 183.405 45.360 183.785 ;
        RECT 46.480 183.405 46.810 183.785 ;
        RECT 47.410 182.945 47.670 183.785 ;
        RECT 47.845 183.240 53.190 183.785 ;
        RECT 49.430 182.410 49.770 183.240 ;
        RECT 53.365 182.965 53.625 183.785 ;
        RECT 55.655 183.325 55.985 183.785 ;
        RECT 57.045 183.405 57.375 183.785 ;
        RECT 58.445 183.405 58.775 183.785 ;
        RECT 59.375 182.985 59.615 183.785 ;
        RECT 59.805 183.015 63.315 183.785 ;
        RECT 64.225 183.250 64.735 183.785 ;
        RECT 66.695 183.385 67.025 183.785 ;
        RECT 67.625 183.060 67.915 183.785 ;
        RECT 69.745 183.250 70.255 183.785 ;
        RECT 72.215 183.385 72.545 183.785 ;
        RECT 73.885 183.250 74.395 183.785 ;
        RECT 76.355 183.385 76.685 183.785 ;
        RECT 77.715 183.385 78.100 183.785 ;
        RECT 79.130 183.385 79.515 183.785 ;
        RECT 80.725 183.385 81.110 183.785 ;
        RECT 82.315 183.385 82.645 183.785 ;
        RECT 84.605 183.250 85.115 183.785 ;
        RECT 86.025 183.015 87.695 183.785 ;
        RECT 88.295 183.385 88.625 183.785 ;
        RECT 90.585 183.250 91.095 183.785 ;
        RECT 92.445 183.405 92.775 183.785 ;
        RECT 93.385 183.060 93.675 183.785 ;
        RECT 94.275 183.385 94.605 183.785 ;
        RECT 96.565 183.250 97.075 183.785 ;
        RECT 98.415 183.385 98.745 183.785 ;
        RECT 100.705 183.250 101.215 183.785 ;
        RECT 59.805 182.495 61.455 183.015 ;
        RECT 86.025 182.495 86.775 183.015 ;
        RECT 102.595 182.985 102.925 183.785 ;
        RECT 103.435 183.305 103.765 183.785 ;
        RECT 104.275 183.305 104.605 183.785 ;
        RECT 105.195 183.305 105.365 183.785 ;
        RECT 106.035 183.305 106.205 183.785 ;
        RECT 107.155 183.385 107.485 183.785 ;
        RECT 109.445 183.250 109.955 183.785 ;
        RECT 111.305 183.305 111.545 183.785 ;
        RECT 112.135 183.305 112.465 183.785 ;
        RECT 112.975 182.985 113.305 183.785 ;
        RECT 114.545 183.035 115.755 183.785 ;
        RECT 115.235 182.495 115.755 183.035 ;
        RECT 41.865 179.265 42.385 179.805 ;
        RECT 41.865 178.515 43.075 179.265 ;
        RECT 44.830 179.060 45.170 179.890 ;
        RECT 43.245 178.515 48.590 179.060 ;
        RECT 50.310 178.515 50.480 179.255 ;
        RECT 52.370 178.515 52.540 178.985 ;
        RECT 53.425 178.515 53.635 179.335 ;
        RECT 54.305 178.515 54.535 179.335 ;
        RECT 54.745 178.515 55.035 179.240 ;
        RECT 56.790 179.060 57.130 179.890 ;
        RECT 60.725 179.285 61.475 179.805 ;
        RECT 55.205 178.515 60.550 179.060 ;
        RECT 60.725 178.515 62.395 179.285 ;
        RECT 69.465 179.265 69.985 179.805 ;
        RECT 73.145 179.285 73.895 179.805 ;
        RECT 76.825 179.285 78.475 179.805 ;
        RECT 63.455 178.515 63.785 178.915 ;
        RECT 65.745 178.515 66.255 179.050 ;
        RECT 68.525 178.515 68.855 178.895 ;
        RECT 69.465 178.515 70.675 179.265 ;
        RECT 70.905 178.515 71.155 178.980 ;
        RECT 71.825 178.515 71.995 178.975 ;
        RECT 72.665 178.515 72.930 178.975 ;
        RECT 73.145 178.515 74.815 179.285 ;
        RECT 74.990 178.515 75.325 178.915 ;
        RECT 75.910 178.515 76.185 178.995 ;
        RECT 76.825 178.515 80.335 179.285 ;
        RECT 80.505 178.515 80.795 179.240 ;
        RECT 82.550 179.060 82.890 179.890 ;
        RECT 86.485 179.285 87.235 179.805 ;
        RECT 80.965 178.515 86.310 179.060 ;
        RECT 86.485 178.515 88.155 179.285 ;
        RECT 89.525 178.515 90.035 179.050 ;
        RECT 91.995 178.515 92.325 178.915 ;
        RECT 93.365 178.515 93.695 178.895 ;
        RECT 95.230 178.515 95.490 179.355 ;
        RECT 115.235 179.265 115.755 179.805 ;
        RECT 96.090 178.515 96.420 178.895 ;
        RECT 97.505 178.515 97.835 178.895 ;
        RECT 98.885 178.515 99.215 178.895 ;
        RECT 100.715 178.515 101.045 178.915 ;
        RECT 103.005 178.515 103.515 179.050 ;
        RECT 104.865 178.515 105.195 178.895 ;
        RECT 106.265 178.515 106.555 179.240 ;
        RECT 107.195 178.515 107.470 178.995 ;
        RECT 108.055 178.515 108.390 178.915 ;
        RECT 109.630 178.515 110.015 178.915 ;
        RECT 111.225 178.515 111.610 178.915 ;
        RECT 112.640 178.515 113.025 178.915 ;
        RECT 114.545 178.515 115.755 179.265 ;
        RECT 41.780 178.345 115.840 178.515 ;
        RECT 41.865 177.595 43.075 178.345 ;
        RECT 43.245 177.800 48.590 178.345 ;
        RECT 50.195 177.885 50.365 178.345 ;
        RECT 51.595 177.885 51.765 178.345 ;
        RECT 52.445 177.800 57.790 178.345 ;
        RECT 58.855 177.945 59.185 178.345 ;
        RECT 61.145 177.810 61.655 178.345 ;
        RECT 63.035 177.865 63.310 178.345 ;
        RECT 63.955 177.865 64.210 178.345 ;
        RECT 64.815 177.865 65.095 178.345 ;
        RECT 41.865 177.055 42.385 177.595 ;
        RECT 44.830 176.970 45.170 177.800 ;
        RECT 54.030 176.970 54.370 177.800 ;
        RECT 65.325 177.575 66.995 178.345 ;
        RECT 67.625 177.620 67.915 178.345 ;
        RECT 69.535 177.885 69.705 178.345 ;
        RECT 70.385 177.800 75.730 178.345 ;
        RECT 76.335 177.945 76.665 178.345 ;
        RECT 78.625 177.810 79.135 178.345 ;
        RECT 80.555 177.885 80.725 178.345 ;
        RECT 83.280 177.965 83.610 178.345 ;
        RECT 84.300 177.885 84.470 178.345 ;
        RECT 65.325 177.055 66.075 177.575 ;
        RECT 71.970 176.970 72.310 177.800 ;
        RECT 86.530 177.625 86.820 178.345 ;
        RECT 88.775 177.965 89.105 178.345 ;
        RECT 90.435 177.885 90.685 178.345 ;
        RECT 92.005 177.595 93.215 178.345 ;
        RECT 93.385 177.620 93.675 178.345 ;
        RECT 94.275 177.945 94.605 178.345 ;
        RECT 96.565 177.810 97.075 178.345 ;
        RECT 98.335 177.865 98.505 178.345 ;
        RECT 99.175 177.865 99.345 178.345 ;
        RECT 99.935 177.865 100.265 178.345 ;
        RECT 100.775 177.865 101.105 178.345 ;
        RECT 92.005 177.055 92.525 177.595 ;
        RECT 101.615 177.545 101.945 178.345 ;
        RECT 103.475 177.945 103.805 178.345 ;
        RECT 105.765 177.810 106.275 178.345 ;
        RECT 107.650 177.505 107.910 178.345 ;
        RECT 108.510 177.965 108.840 178.345 ;
        RECT 110.415 177.545 110.745 178.345 ;
        RECT 111.255 177.865 111.585 178.345 ;
        RECT 112.095 177.865 112.425 178.345 ;
        RECT 113.015 177.865 113.185 178.345 ;
        RECT 113.855 177.865 114.025 178.345 ;
        RECT 114.545 177.595 115.755 178.345 ;
        RECT 115.235 177.055 115.755 177.595 ;
        RECT 41.865 173.825 42.385 174.365 ;
        RECT 41.865 173.075 43.075 173.825 ;
        RECT 44.830 173.620 45.170 174.450 ;
        RECT 43.245 173.075 48.590 173.620 ;
        RECT 49.735 173.075 49.905 173.895 ;
        RECT 51.985 173.845 53.195 174.365 ;
        RECT 50.575 173.075 50.925 173.465 ;
        RECT 51.985 173.075 54.575 173.845 ;
        RECT 54.745 173.075 55.035 173.800 ;
        RECT 56.175 173.075 56.345 173.895 ;
        RECT 60.725 173.825 61.245 174.365 ;
        RECT 86.485 173.845 87.235 174.365 ;
        RECT 57.015 173.075 57.365 173.465 ;
        RECT 59.155 173.075 59.405 173.535 ;
        RECT 60.725 173.075 61.935 173.825 ;
        RECT 62.845 173.075 63.355 173.610 ;
        RECT 65.315 173.075 65.645 173.475 ;
        RECT 66.675 173.075 67.005 173.475 ;
        RECT 68.965 173.075 69.475 173.610 ;
        RECT 70.815 173.075 71.145 173.455 ;
        RECT 73.100 173.075 73.390 173.795 ;
        RECT 75.450 173.075 75.620 173.535 ;
        RECT 76.310 173.075 76.640 173.455 ;
        RECT 79.195 173.075 79.365 173.535 ;
        RECT 80.505 173.075 80.795 173.800 ;
        RECT 81.705 173.075 82.215 173.610 ;
        RECT 84.175 173.075 84.505 173.475 ;
        RECT 85.545 173.075 85.875 173.455 ;
        RECT 86.485 173.075 88.155 173.845 ;
        RECT 89.065 173.075 89.575 173.610 ;
        RECT 91.535 173.075 91.865 173.475 ;
        RECT 93.205 173.075 93.715 173.610 ;
        RECT 95.675 173.075 96.005 173.475 ;
        RECT 97.955 173.075 98.285 173.475 ;
        RECT 100.245 173.075 100.755 173.610 ;
        RECT 102.095 173.075 102.425 173.475 ;
        RECT 104.385 173.075 104.895 173.610 ;
        RECT 106.265 173.075 106.555 173.800 ;
        RECT 107.155 173.075 107.485 173.475 ;
        RECT 109.445 173.075 109.955 173.610 ;
        RECT 111.935 173.075 112.265 173.875 ;
        RECT 115.235 173.825 115.755 174.365 ;
        RECT 112.775 173.075 113.105 173.555 ;
        RECT 113.695 173.075 113.935 173.555 ;
        RECT 114.545 173.075 115.755 173.825 ;
        RECT 41.780 172.905 115.840 173.075 ;
        RECT 41.865 172.155 43.075 172.905 ;
        RECT 43.245 172.360 48.590 172.905 ;
        RECT 48.765 172.360 54.110 172.905 ;
        RECT 41.865 171.615 42.385 172.155 ;
        RECT 44.830 171.530 45.170 172.360 ;
        RECT 50.350 171.530 50.690 172.360 ;
        RECT 54.285 172.135 55.955 172.905 ;
        RECT 56.555 172.505 56.885 172.905 ;
        RECT 58.845 172.370 59.355 172.905 ;
        RECT 60.265 172.135 61.935 172.905 ;
        RECT 63.355 172.505 63.685 172.905 ;
        RECT 65.025 172.520 65.360 172.905 ;
        RECT 66.245 172.155 67.455 172.905 ;
        RECT 67.625 172.180 67.915 172.905 ;
        RECT 68.525 172.525 68.855 172.905 ;
        RECT 69.465 172.360 74.810 172.905 ;
        RECT 74.985 172.360 80.330 172.905 ;
        RECT 81.395 172.505 81.725 172.905 ;
        RECT 83.685 172.370 84.195 172.905 ;
        RECT 87.060 172.500 87.390 172.905 ;
        RECT 88.800 172.445 89.145 172.905 ;
        RECT 89.815 172.445 89.985 172.905 ;
        RECT 90.655 172.445 90.825 172.905 ;
        RECT 54.285 171.615 55.035 172.135 ;
        RECT 60.265 171.615 61.015 172.135 ;
        RECT 66.245 171.615 66.765 172.155 ;
        RECT 71.050 171.530 71.390 172.360 ;
        RECT 76.570 171.530 76.910 172.360 ;
        RECT 91.085 172.135 92.755 172.905 ;
        RECT 93.385 172.180 93.675 172.905 ;
        RECT 93.845 172.135 96.435 172.905 ;
        RECT 98.100 172.500 98.430 172.905 ;
        RECT 99.840 172.445 100.185 172.905 ;
        RECT 100.855 172.445 101.025 172.905 ;
        RECT 101.695 172.445 101.865 172.905 ;
        RECT 102.125 172.135 104.715 172.905 ;
        RECT 105.315 172.525 105.645 172.905 ;
        RECT 107.600 172.185 107.890 172.905 ;
        RECT 109.950 172.445 110.120 172.905 ;
        RECT 110.810 172.525 111.140 172.905 ;
        RECT 113.695 172.445 113.865 172.905 ;
        RECT 114.545 172.155 115.755 172.905 ;
        RECT 91.085 171.615 91.835 172.135 ;
        RECT 93.845 171.615 95.055 172.135 ;
        RECT 102.125 171.615 103.335 172.135 ;
        RECT 115.235 171.615 115.755 172.155 ;
        RECT 41.865 168.385 42.385 168.925 ;
        RECT 41.865 167.635 43.075 168.385 ;
        RECT 44.830 168.180 45.170 169.010 ;
        RECT 50.350 168.180 50.690 169.010 ;
        RECT 55.205 168.405 56.855 168.925 ;
        RECT 43.245 167.635 48.590 168.180 ;
        RECT 48.765 167.635 54.110 168.180 ;
        RECT 54.745 167.635 55.035 168.360 ;
        RECT 55.205 167.635 58.715 168.405 ;
        RECT 58.885 168.385 59.405 168.925 ;
        RECT 64.405 168.405 65.615 168.925 ;
        RECT 58.885 167.635 60.095 168.385 ;
        RECT 61.005 167.635 61.515 168.170 ;
        RECT 63.475 167.635 63.805 168.035 ;
        RECT 64.405 167.635 66.995 168.405 ;
        RECT 68.515 167.635 68.845 168.035 ;
        RECT 70.175 167.635 70.505 168.035 ;
        RECT 71.325 167.635 71.595 168.455 ;
        RECT 75.905 168.405 77.555 168.925 ;
        RECT 72.195 167.635 72.525 168.035 ;
        RECT 74.485 167.635 74.995 168.170 ;
        RECT 75.905 167.635 79.415 168.405 ;
        RECT 80.505 167.635 80.795 168.360 ;
        RECT 82.315 167.635 82.645 168.015 ;
        RECT 84.600 167.635 84.890 168.355 ;
        RECT 86.950 167.635 87.120 168.095 ;
        RECT 87.810 167.635 88.140 168.015 ;
        RECT 90.695 167.635 90.865 168.095 ;
        RECT 93.355 167.635 93.685 168.035 ;
        RECT 95.015 167.635 95.345 168.035 ;
        RECT 96.165 167.635 96.435 168.455 ;
        RECT 115.235 168.385 115.755 168.925 ;
        RECT 97.035 167.635 97.365 168.015 ;
        RECT 99.320 167.635 99.610 168.355 ;
        RECT 101.670 167.635 101.840 168.095 ;
        RECT 102.530 167.635 102.860 168.015 ;
        RECT 105.415 167.635 105.585 168.095 ;
        RECT 106.265 167.635 106.555 168.360 ;
        RECT 107.155 167.635 107.485 168.035 ;
        RECT 109.445 167.635 109.955 168.170 ;
        RECT 111.305 167.635 111.635 168.015 ;
        RECT 112.685 167.635 113.015 168.015 ;
        RECT 114.545 167.635 115.755 168.385 ;
        RECT 41.780 167.465 115.840 167.635 ;
        RECT 41.865 166.715 43.075 167.465 ;
        RECT 43.245 166.920 48.590 167.465 ;
        RECT 41.865 166.175 42.385 166.715 ;
        RECT 44.830 166.090 45.170 166.920 ;
        RECT 48.765 166.695 50.435 167.465 ;
        RECT 51.115 167.005 51.285 167.465 ;
        RECT 53.840 167.085 54.170 167.465 ;
        RECT 54.860 167.005 55.030 167.465 ;
        RECT 57.090 166.745 57.380 167.465 ;
        RECT 59.335 167.085 59.665 167.465 ;
        RECT 60.265 166.920 65.610 167.465 ;
        RECT 48.765 166.175 49.515 166.695 ;
        RECT 61.850 166.090 62.190 166.920 ;
        RECT 65.785 166.695 67.455 167.465 ;
        RECT 67.625 166.740 67.915 167.465 ;
        RECT 68.085 166.695 70.675 167.465 ;
        RECT 70.850 167.065 71.185 167.465 ;
        RECT 71.770 166.985 72.045 167.465 ;
        RECT 72.685 166.695 74.355 167.465 ;
        RECT 75.315 167.065 75.645 167.465 ;
        RECT 76.985 167.080 77.320 167.465 ;
        RECT 78.205 166.715 79.415 167.465 ;
        RECT 79.590 167.065 79.925 167.465 ;
        RECT 80.510 166.985 80.785 167.465 ;
        RECT 81.425 166.920 86.770 167.465 ;
        RECT 65.785 166.175 66.535 166.695 ;
        RECT 68.085 166.175 69.295 166.695 ;
        RECT 72.685 166.175 73.435 166.695 ;
        RECT 78.205 166.175 78.725 166.715 ;
        RECT 83.010 166.090 83.350 166.920 ;
        RECT 86.945 166.695 90.455 167.465 ;
        RECT 91.550 167.065 91.885 167.465 ;
        RECT 92.470 166.985 92.745 167.465 ;
        RECT 93.385 166.740 93.675 167.465 ;
        RECT 94.735 167.065 95.065 167.465 ;
        RECT 96.395 167.065 96.725 167.465 ;
        RECT 86.945 166.175 88.595 166.695 ;
        RECT 97.545 166.645 97.815 167.465 ;
        RECT 97.985 166.920 103.330 167.465 ;
        RECT 104.515 167.005 104.685 167.465 ;
        RECT 105.355 167.005 105.525 167.465 ;
        RECT 106.195 167.005 106.540 167.465 ;
        RECT 107.950 167.060 108.280 167.465 ;
        RECT 110.375 167.065 110.705 167.465 ;
        RECT 112.665 166.930 113.175 167.465 ;
        RECT 99.570 166.090 99.910 166.920 ;
        RECT 114.545 166.715 115.755 167.465 ;
        RECT 115.235 166.175 115.755 166.715 ;
        RECT 41.865 162.945 42.385 163.485 ;
        RECT 41.865 162.195 43.075 162.945 ;
        RECT 44.830 162.740 45.170 163.570 ;
        RECT 50.350 162.740 50.690 163.570 ;
        RECT 43.245 162.195 48.590 162.740 ;
        RECT 48.765 162.195 54.110 162.740 ;
        RECT 54.745 162.195 55.035 162.920 ;
        RECT 56.095 162.195 56.445 162.585 ;
        RECT 57.115 162.195 57.285 163.015 ;
        RECT 58.425 162.965 59.635 163.485 ;
        RECT 58.425 162.195 61.015 162.965 ;
        RECT 61.695 162.195 61.865 162.655 ;
        RECT 64.420 162.195 64.750 162.575 ;
        RECT 65.440 162.195 65.610 162.655 ;
        RECT 67.670 162.195 67.960 162.915 ;
        RECT 72.430 162.740 72.770 163.570 ;
        RECT 76.365 162.965 77.115 163.485 ;
        RECT 69.915 162.195 70.245 162.575 ;
        RECT 70.845 162.195 76.190 162.740 ;
        RECT 76.365 162.195 78.035 162.965 ;
        RECT 78.670 162.195 79.005 162.595 ;
        RECT 79.590 162.195 79.865 162.675 ;
        RECT 80.505 162.195 80.795 162.920 ;
        RECT 81.855 162.195 82.185 162.595 ;
        RECT 83.515 162.195 83.845 162.595 ;
        RECT 84.665 162.195 84.935 163.015 ;
        RECT 90.165 162.965 91.815 163.485 ;
        RECT 103.965 162.965 104.715 163.485 ;
        RECT 106.725 162.965 107.935 163.485 ;
        RECT 86.455 162.195 86.785 162.595 ;
        RECT 88.745 162.195 89.255 162.730 ;
        RECT 90.165 162.195 93.675 162.965 ;
        RECT 94.275 162.195 94.605 162.595 ;
        RECT 96.565 162.195 97.075 162.730 ;
        RECT 98.415 162.195 98.745 162.595 ;
        RECT 100.705 162.195 101.215 162.730 ;
        RECT 102.595 162.195 102.870 162.675 ;
        RECT 103.455 162.195 103.790 162.595 ;
        RECT 103.965 162.195 105.635 162.965 ;
        RECT 106.265 162.195 106.555 162.920 ;
        RECT 106.725 162.195 109.315 162.965 ;
        RECT 115.235 162.945 115.755 163.485 ;
        RECT 109.925 162.195 110.255 162.575 ;
        RECT 111.305 162.195 111.635 162.575 ;
        RECT 112.685 162.195 113.015 162.575 ;
        RECT 114.545 162.195 115.755 162.945 ;
        RECT 41.780 162.025 115.840 162.195 ;
        RECT 41.865 161.275 43.075 162.025 ;
        RECT 43.245 161.480 48.590 162.025 ;
        RECT 41.865 160.735 42.385 161.275 ;
        RECT 44.830 160.650 45.170 161.480 ;
        RECT 48.765 161.255 51.355 162.025 ;
        RECT 52.035 161.635 52.365 162.025 ;
        RECT 52.875 161.635 53.205 162.025 ;
        RECT 48.765 160.735 49.975 161.255 ;
        RECT 54.745 161.190 55.035 162.025 ;
        RECT 56.175 161.205 56.345 162.025 ;
        RECT 57.015 161.635 57.365 162.025 ;
        RECT 58.425 161.255 61.015 162.025 ;
        RECT 58.425 160.735 59.635 161.255 ;
        RECT 62.155 161.205 62.325 162.025 ;
        RECT 62.995 161.635 63.345 162.025 ;
        RECT 64.455 161.635 64.785 162.025 ;
        RECT 65.295 161.635 65.625 162.025 ;
        RECT 67.165 161.190 67.455 162.025 ;
        RECT 67.625 161.300 67.915 162.025 ;
        RECT 68.085 161.255 69.755 162.025 ;
        RECT 70.355 161.625 70.685 162.025 ;
        RECT 72.645 161.490 73.155 162.025 ;
        RECT 74.495 161.625 74.825 162.025 ;
        RECT 76.785 161.490 77.295 162.025 ;
        RECT 68.085 160.735 68.835 161.255 ;
        RECT 80.095 161.205 80.265 162.025 ;
        RECT 80.935 161.635 81.285 162.025 ;
        RECT 82.345 161.480 87.690 162.025 ;
        RECT 83.930 160.650 84.270 161.480 ;
        RECT 87.865 161.255 89.535 162.025 ;
        RECT 87.865 160.735 88.615 161.255 ;
        RECT 89.705 161.190 89.995 162.025 ;
        RECT 91.535 161.635 91.865 162.025 ;
        RECT 92.375 161.635 92.705 162.025 ;
        RECT 93.385 161.300 93.675 162.025 ;
        RECT 93.845 161.255 95.515 162.025 ;
        RECT 95.690 161.625 96.025 162.025 ;
        RECT 96.610 161.545 96.885 162.025 ;
        RECT 97.525 161.255 101.035 162.025 ;
        RECT 102.095 161.625 102.425 162.025 ;
        RECT 104.385 161.490 104.895 162.025 ;
        RECT 106.520 161.640 106.855 162.025 ;
        RECT 108.195 161.625 108.525 162.025 ;
        RECT 109.485 161.275 110.695 162.025 ;
        RECT 111.305 161.645 111.635 162.025 ;
        RECT 112.685 161.645 113.015 162.025 ;
        RECT 114.545 161.275 115.755 162.025 ;
        RECT 93.845 160.735 94.595 161.255 ;
        RECT 97.525 160.735 99.175 161.255 ;
        RECT 109.485 160.735 110.005 161.275 ;
        RECT 115.235 160.735 115.755 161.275 ;
        RECT 41.865 157.505 42.385 158.045 ;
        RECT 45.085 157.525 46.735 158.045 ;
        RECT 50.145 157.525 51.795 158.045 ;
        RECT 56.585 157.525 57.335 158.045 ;
        RECT 60.265 157.525 61.915 158.045 ;
        RECT 65.325 157.525 66.075 158.045 ;
        RECT 41.865 156.755 43.075 157.505 ;
        RECT 44.145 156.755 44.475 157.135 ;
        RECT 45.085 156.755 48.595 157.525 ;
        RECT 49.205 156.755 49.535 157.135 ;
        RECT 50.145 156.755 53.655 157.525 ;
        RECT 54.745 156.755 55.035 157.480 ;
        RECT 55.645 156.755 55.975 157.135 ;
        RECT 56.585 156.755 58.255 157.525 ;
        RECT 59.325 156.755 59.655 157.135 ;
        RECT 60.265 156.755 63.775 157.525 ;
        RECT 64.385 156.755 64.715 157.135 ;
        RECT 65.325 156.755 66.995 157.525 ;
        RECT 67.625 156.755 67.915 157.480 ;
        RECT 69.055 156.755 69.225 157.575 ;
        RECT 72.685 157.505 73.205 158.045 ;
        RECT 75.445 157.525 77.095 158.045 ;
        RECT 80.965 157.525 81.715 158.045 ;
        RECT 69.895 156.755 70.245 157.145 ;
        RECT 71.745 156.755 72.075 157.135 ;
        RECT 72.685 156.755 73.895 157.505 ;
        RECT 74.505 156.755 74.835 157.135 ;
        RECT 75.445 156.755 78.955 157.525 ;
        RECT 79.565 156.755 79.895 157.135 ;
        RECT 80.505 156.755 80.795 157.480 ;
        RECT 80.965 156.755 82.635 157.525 ;
        RECT 84.155 156.755 84.505 157.145 ;
        RECT 85.175 156.755 85.345 157.575 ;
        RECT 87.865 157.505 88.385 158.045 ;
        RECT 90.625 157.525 91.835 158.045 ;
        RECT 95.685 157.525 97.335 158.045 ;
        RECT 100.745 157.525 102.395 158.045 ;
        RECT 86.925 156.755 87.255 157.135 ;
        RECT 87.865 156.755 89.075 157.505 ;
        RECT 89.685 156.755 90.015 157.135 ;
        RECT 90.625 156.755 93.215 157.525 ;
        RECT 93.385 156.755 93.675 157.480 ;
        RECT 94.745 156.755 95.075 157.135 ;
        RECT 95.685 156.755 99.195 157.525 ;
        RECT 99.805 156.755 100.135 157.135 ;
        RECT 100.745 156.755 104.255 157.525 ;
        RECT 104.865 156.755 105.195 157.135 ;
        RECT 106.265 156.755 106.555 157.480 ;
        RECT 107.615 156.755 107.945 157.155 ;
        RECT 109.275 156.755 109.605 157.155 ;
        RECT 110.425 156.755 110.695 157.575 ;
        RECT 115.235 157.505 115.755 158.045 ;
        RECT 111.305 156.755 111.635 157.135 ;
        RECT 113.605 156.755 113.935 157.135 ;
        RECT 114.545 156.755 115.755 157.505 ;
        RECT 41.780 156.585 115.840 156.755 ;
        RECT 63.940 125.510 64.110 127.550 ;
        RECT 64.530 125.510 64.700 127.550 ;
        RECT 70.170 125.510 70.340 127.550 ;
        RECT 72.050 125.510 72.220 127.550 ;
        RECT 73.930 125.510 74.100 127.550 ;
        RECT 76.650 126.690 76.860 127.060 ;
        RECT 76.650 125.400 76.860 125.770 ;
        RECT 86.600 125.510 86.770 127.550 ;
        RECT 87.190 125.510 87.360 127.550 ;
        RECT 92.830 125.510 93.000 127.550 ;
        RECT 94.710 125.510 94.880 127.550 ;
        RECT 96.590 125.510 96.760 127.550 ;
        RECT 99.310 126.690 99.520 127.060 ;
        RECT 99.310 125.400 99.520 125.770 ;
        RECT 109.260 125.510 109.430 127.550 ;
        RECT 109.850 125.510 110.020 127.550 ;
        RECT 115.490 125.510 115.660 127.550 ;
        RECT 117.370 125.510 117.540 127.550 ;
        RECT 119.250 125.510 119.420 127.550 ;
        RECT 121.970 126.690 122.180 127.060 ;
        RECT 121.970 125.400 122.180 125.770 ;
        RECT 124.200 124.620 124.550 126.780 ;
        RECT 58.060 122.525 58.430 122.735 ;
        RECT 63.940 122.420 64.110 124.460 ;
        RECT 64.530 122.420 64.700 124.460 ;
        RECT 70.170 122.420 70.340 124.460 ;
        RECT 72.050 122.420 72.220 124.460 ;
        RECT 73.930 122.420 74.100 124.460 ;
        RECT 76.650 124.115 76.860 124.485 ;
        RECT 76.650 122.830 76.860 123.200 ;
        RECT 80.720 122.525 81.090 122.735 ;
        RECT 86.600 122.420 86.770 124.460 ;
        RECT 87.190 122.420 87.360 124.460 ;
        RECT 92.830 122.420 93.000 124.460 ;
        RECT 94.710 122.420 94.880 124.460 ;
        RECT 96.590 122.420 96.760 124.460 ;
        RECT 99.310 124.115 99.520 124.485 ;
        RECT 99.310 122.830 99.520 123.200 ;
        RECT 103.380 122.525 103.750 122.735 ;
        RECT 109.260 122.420 109.430 124.460 ;
        RECT 109.850 122.420 110.020 124.460 ;
        RECT 115.490 122.420 115.660 124.460 ;
        RECT 117.370 122.420 117.540 124.460 ;
        RECT 119.250 122.420 119.420 124.460 ;
        RECT 121.970 124.115 122.180 124.485 ;
        RECT 121.970 122.830 122.180 123.200 ;
        RECT 59.470 121.620 59.640 122.160 ;
        RECT 60.870 121.620 61.040 122.160 ;
        RECT 82.130 121.620 82.300 122.160 ;
        RECT 83.530 121.620 83.700 122.160 ;
        RECT 104.790 121.620 104.960 122.160 ;
        RECT 106.190 121.620 106.360 122.160 ;
        RECT 41.280 108.170 41.450 110.210 ;
        RECT 41.870 108.170 42.040 110.210 ;
        RECT 47.510 108.170 47.680 110.210 ;
        RECT 49.390 108.170 49.560 110.210 ;
        RECT 51.270 108.170 51.440 110.210 ;
        RECT 53.990 109.350 54.200 109.720 ;
        RECT 53.990 108.060 54.200 108.430 ;
        RECT 63.940 108.170 64.110 110.210 ;
        RECT 64.530 108.170 64.700 110.210 ;
        RECT 70.170 108.170 70.340 110.210 ;
        RECT 72.050 108.170 72.220 110.210 ;
        RECT 73.930 108.170 74.100 110.210 ;
        RECT 76.650 109.350 76.860 109.720 ;
        RECT 76.650 108.060 76.860 108.430 ;
        RECT 86.600 108.170 86.770 110.210 ;
        RECT 87.190 108.170 87.360 110.210 ;
        RECT 92.830 108.170 93.000 110.210 ;
        RECT 94.710 108.170 94.880 110.210 ;
        RECT 96.590 108.170 96.760 110.210 ;
        RECT 99.310 109.350 99.520 109.720 ;
        RECT 99.310 108.060 99.520 108.430 ;
        RECT 109.260 108.170 109.430 110.210 ;
        RECT 109.850 108.170 110.020 110.210 ;
        RECT 115.490 108.170 115.660 110.210 ;
        RECT 117.370 108.170 117.540 110.210 ;
        RECT 119.250 108.170 119.420 110.210 ;
        RECT 121.970 109.350 122.180 109.720 ;
        RECT 121.970 108.060 122.180 108.430 ;
        RECT 35.400 105.185 35.770 105.395 ;
        RECT 41.280 105.080 41.450 107.120 ;
        RECT 41.870 105.080 42.040 107.120 ;
        RECT 47.510 105.080 47.680 107.120 ;
        RECT 49.390 105.080 49.560 107.120 ;
        RECT 51.270 105.080 51.440 107.120 ;
        RECT 53.990 106.775 54.200 107.145 ;
        RECT 53.990 105.490 54.200 105.860 ;
        RECT 58.060 105.185 58.430 105.395 ;
        RECT 63.940 105.080 64.110 107.120 ;
        RECT 64.530 105.080 64.700 107.120 ;
        RECT 70.170 105.080 70.340 107.120 ;
        RECT 72.050 105.080 72.220 107.120 ;
        RECT 73.930 105.080 74.100 107.120 ;
        RECT 76.650 106.775 76.860 107.145 ;
        RECT 76.650 105.490 76.860 105.860 ;
        RECT 80.720 105.185 81.090 105.395 ;
        RECT 86.600 105.080 86.770 107.120 ;
        RECT 87.190 105.080 87.360 107.120 ;
        RECT 92.830 105.080 93.000 107.120 ;
        RECT 94.710 105.080 94.880 107.120 ;
        RECT 96.590 105.080 96.760 107.120 ;
        RECT 99.310 106.775 99.520 107.145 ;
        RECT 99.310 105.490 99.520 105.860 ;
        RECT 103.380 105.185 103.750 105.395 ;
        RECT 109.260 105.080 109.430 107.120 ;
        RECT 109.850 105.080 110.020 107.120 ;
        RECT 115.490 105.080 115.660 107.120 ;
        RECT 117.370 105.080 117.540 107.120 ;
        RECT 119.250 105.080 119.420 107.120 ;
        RECT 121.970 106.775 122.180 107.145 ;
        RECT 121.970 105.490 122.180 105.860 ;
        RECT 36.810 104.280 36.980 104.820 ;
        RECT 38.210 104.280 38.380 104.820 ;
        RECT 59.470 104.280 59.640 104.820 ;
        RECT 60.870 104.280 61.040 104.820 ;
        RECT 82.130 104.280 82.300 104.820 ;
        RECT 83.530 104.280 83.700 104.820 ;
        RECT 104.790 104.280 104.960 104.820 ;
        RECT 106.190 104.280 106.360 104.820 ;
        RECT 41.280 90.830 41.450 92.870 ;
        RECT 41.870 90.830 42.040 92.870 ;
        RECT 47.510 90.830 47.680 92.870 ;
        RECT 49.390 90.830 49.560 92.870 ;
        RECT 51.270 90.830 51.440 92.870 ;
        RECT 53.990 92.010 54.200 92.380 ;
        RECT 53.990 90.720 54.200 91.090 ;
        RECT 63.940 90.830 64.110 92.870 ;
        RECT 64.530 90.830 64.700 92.870 ;
        RECT 70.170 90.830 70.340 92.870 ;
        RECT 72.050 90.830 72.220 92.870 ;
        RECT 73.930 90.830 74.100 92.870 ;
        RECT 76.650 92.010 76.860 92.380 ;
        RECT 76.650 90.720 76.860 91.090 ;
        RECT 86.600 90.830 86.770 92.870 ;
        RECT 87.190 90.830 87.360 92.870 ;
        RECT 92.830 90.830 93.000 92.870 ;
        RECT 94.710 90.830 94.880 92.870 ;
        RECT 96.590 90.830 96.760 92.870 ;
        RECT 99.310 92.010 99.520 92.380 ;
        RECT 99.310 90.720 99.520 91.090 ;
        RECT 109.260 90.830 109.430 92.870 ;
        RECT 109.850 90.830 110.020 92.870 ;
        RECT 115.490 90.830 115.660 92.870 ;
        RECT 117.370 90.830 117.540 92.870 ;
        RECT 119.250 90.830 119.420 92.870 ;
        RECT 121.970 92.010 122.180 92.380 ;
        RECT 121.970 90.720 122.180 91.090 ;
        RECT 35.400 87.845 35.770 88.055 ;
        RECT 41.280 87.740 41.450 89.780 ;
        RECT 41.870 87.740 42.040 89.780 ;
        RECT 47.510 87.740 47.680 89.780 ;
        RECT 49.390 87.740 49.560 89.780 ;
        RECT 51.270 87.740 51.440 89.780 ;
        RECT 53.990 89.435 54.200 89.805 ;
        RECT 53.990 88.150 54.200 88.520 ;
        RECT 58.060 87.845 58.430 88.055 ;
        RECT 63.940 87.740 64.110 89.780 ;
        RECT 64.530 87.740 64.700 89.780 ;
        RECT 70.170 87.740 70.340 89.780 ;
        RECT 72.050 87.740 72.220 89.780 ;
        RECT 73.930 87.740 74.100 89.780 ;
        RECT 76.650 89.435 76.860 89.805 ;
        RECT 76.650 88.150 76.860 88.520 ;
        RECT 80.720 87.845 81.090 88.055 ;
        RECT 86.600 87.740 86.770 89.780 ;
        RECT 87.190 87.740 87.360 89.780 ;
        RECT 92.830 87.740 93.000 89.780 ;
        RECT 94.710 87.740 94.880 89.780 ;
        RECT 96.590 87.740 96.760 89.780 ;
        RECT 99.310 89.435 99.520 89.805 ;
        RECT 99.310 88.150 99.520 88.520 ;
        RECT 103.380 87.845 103.750 88.055 ;
        RECT 109.260 87.740 109.430 89.780 ;
        RECT 109.850 87.740 110.020 89.780 ;
        RECT 115.490 87.740 115.660 89.780 ;
        RECT 117.370 87.740 117.540 89.780 ;
        RECT 119.250 87.740 119.420 89.780 ;
        RECT 121.970 89.435 122.180 89.805 ;
        RECT 121.970 88.150 122.180 88.520 ;
        RECT 36.810 86.940 36.980 87.480 ;
        RECT 38.210 86.940 38.380 87.480 ;
        RECT 59.470 86.940 59.640 87.480 ;
        RECT 60.870 86.940 61.040 87.480 ;
        RECT 82.130 86.940 82.300 87.480 ;
        RECT 83.530 86.940 83.700 87.480 ;
        RECT 104.790 86.940 104.960 87.480 ;
        RECT 106.190 86.940 106.360 87.480 ;
        RECT 41.280 73.490 41.450 75.530 ;
        RECT 41.870 73.490 42.040 75.530 ;
        RECT 47.510 73.490 47.680 75.530 ;
        RECT 49.390 73.490 49.560 75.530 ;
        RECT 51.270 73.490 51.440 75.530 ;
        RECT 53.990 74.670 54.200 75.040 ;
        RECT 53.990 73.380 54.200 73.750 ;
        RECT 63.940 73.490 64.110 75.530 ;
        RECT 64.530 73.490 64.700 75.530 ;
        RECT 70.170 73.490 70.340 75.530 ;
        RECT 72.050 73.490 72.220 75.530 ;
        RECT 73.930 73.490 74.100 75.530 ;
        RECT 76.650 74.670 76.860 75.040 ;
        RECT 76.650 73.380 76.860 73.750 ;
        RECT 86.600 73.490 86.770 75.530 ;
        RECT 87.190 73.490 87.360 75.530 ;
        RECT 92.830 73.490 93.000 75.530 ;
        RECT 94.710 73.490 94.880 75.530 ;
        RECT 96.590 73.490 96.760 75.530 ;
        RECT 99.310 74.670 99.520 75.040 ;
        RECT 99.310 73.380 99.520 73.750 ;
        RECT 109.260 73.490 109.430 75.530 ;
        RECT 109.850 73.490 110.020 75.530 ;
        RECT 115.490 73.490 115.660 75.530 ;
        RECT 117.370 73.490 117.540 75.530 ;
        RECT 119.250 73.490 119.420 75.530 ;
        RECT 121.970 74.670 122.180 75.040 ;
        RECT 121.970 73.380 122.180 73.750 ;
        RECT 35.400 70.505 35.770 70.715 ;
        RECT 41.280 70.400 41.450 72.440 ;
        RECT 41.870 70.400 42.040 72.440 ;
        RECT 47.510 70.400 47.680 72.440 ;
        RECT 49.390 70.400 49.560 72.440 ;
        RECT 51.270 70.400 51.440 72.440 ;
        RECT 53.990 72.095 54.200 72.465 ;
        RECT 53.990 70.810 54.200 71.180 ;
        RECT 58.060 70.505 58.430 70.715 ;
        RECT 63.940 70.400 64.110 72.440 ;
        RECT 64.530 70.400 64.700 72.440 ;
        RECT 70.170 70.400 70.340 72.440 ;
        RECT 72.050 70.400 72.220 72.440 ;
        RECT 73.930 70.400 74.100 72.440 ;
        RECT 76.650 72.095 76.860 72.465 ;
        RECT 76.650 70.810 76.860 71.180 ;
        RECT 80.720 70.505 81.090 70.715 ;
        RECT 86.600 70.400 86.770 72.440 ;
        RECT 87.190 70.400 87.360 72.440 ;
        RECT 92.830 70.400 93.000 72.440 ;
        RECT 94.710 70.400 94.880 72.440 ;
        RECT 96.590 70.400 96.760 72.440 ;
        RECT 99.310 72.095 99.520 72.465 ;
        RECT 99.310 70.810 99.520 71.180 ;
        RECT 103.380 70.505 103.750 70.715 ;
        RECT 109.260 70.400 109.430 72.440 ;
        RECT 109.850 70.400 110.020 72.440 ;
        RECT 115.490 70.400 115.660 72.440 ;
        RECT 117.370 70.400 117.540 72.440 ;
        RECT 119.250 70.400 119.420 72.440 ;
        RECT 121.970 72.095 122.180 72.465 ;
        RECT 121.970 70.810 122.180 71.180 ;
        RECT 36.810 69.600 36.980 70.140 ;
        RECT 38.210 69.600 38.380 70.140 ;
        RECT 59.470 69.600 59.640 70.140 ;
        RECT 60.870 69.600 61.040 70.140 ;
        RECT 82.130 69.600 82.300 70.140 ;
        RECT 83.530 69.600 83.700 70.140 ;
        RECT 104.790 69.600 104.960 70.140 ;
        RECT 106.190 69.600 106.360 70.140 ;
        RECT 41.280 55.490 41.450 57.530 ;
        RECT 41.870 55.490 42.040 57.530 ;
        RECT 47.510 55.490 47.680 57.530 ;
        RECT 49.390 55.490 49.560 57.530 ;
        RECT 51.270 55.490 51.440 57.530 ;
        RECT 53.990 56.670 54.200 57.040 ;
        RECT 53.990 55.380 54.200 55.750 ;
        RECT 63.940 55.490 64.110 57.530 ;
        RECT 64.530 55.490 64.700 57.530 ;
        RECT 70.170 55.490 70.340 57.530 ;
        RECT 72.050 55.490 72.220 57.530 ;
        RECT 73.930 55.490 74.100 57.530 ;
        RECT 76.650 56.670 76.860 57.040 ;
        RECT 76.650 55.380 76.860 55.750 ;
        RECT 86.600 55.490 86.770 57.530 ;
        RECT 87.190 55.490 87.360 57.530 ;
        RECT 92.830 55.490 93.000 57.530 ;
        RECT 94.710 55.490 94.880 57.530 ;
        RECT 96.590 55.490 96.760 57.530 ;
        RECT 99.310 56.670 99.520 57.040 ;
        RECT 99.310 55.380 99.520 55.750 ;
        RECT 109.260 55.490 109.430 57.530 ;
        RECT 109.850 55.490 110.020 57.530 ;
        RECT 115.490 55.490 115.660 57.530 ;
        RECT 117.370 55.490 117.540 57.530 ;
        RECT 119.250 55.490 119.420 57.530 ;
        RECT 121.970 56.670 122.180 57.040 ;
        RECT 121.970 55.380 122.180 55.750 ;
        RECT 41.280 52.400 41.450 54.440 ;
        RECT 41.870 52.400 42.040 54.440 ;
        RECT 47.510 52.400 47.680 54.440 ;
        RECT 49.390 52.400 49.560 54.440 ;
        RECT 51.270 52.400 51.440 54.440 ;
        RECT 53.990 54.095 54.200 54.465 ;
        RECT 53.990 52.810 54.200 53.180 ;
        RECT 63.940 52.400 64.110 54.440 ;
        RECT 64.530 52.400 64.700 54.440 ;
        RECT 70.170 52.400 70.340 54.440 ;
        RECT 72.050 52.400 72.220 54.440 ;
        RECT 73.930 52.400 74.100 54.440 ;
        RECT 76.650 54.095 76.860 54.465 ;
        RECT 76.650 52.810 76.860 53.180 ;
        RECT 86.600 52.400 86.770 54.440 ;
        RECT 87.190 52.400 87.360 54.440 ;
        RECT 92.830 52.400 93.000 54.440 ;
        RECT 94.710 52.400 94.880 54.440 ;
        RECT 96.590 52.400 96.760 54.440 ;
        RECT 99.310 54.095 99.520 54.465 ;
        RECT 99.310 52.810 99.520 53.180 ;
        RECT 109.260 52.400 109.430 54.440 ;
        RECT 109.850 52.400 110.020 54.440 ;
        RECT 115.490 52.400 115.660 54.440 ;
        RECT 117.370 52.400 117.540 54.440 ;
        RECT 119.250 52.400 119.420 54.440 ;
        RECT 121.970 54.095 122.180 54.465 ;
        RECT 121.970 52.810 122.180 53.180 ;
      LAYER mcon ;
        RECT 41.925 183.785 42.095 183.955 ;
        RECT 42.385 183.785 42.555 183.955 ;
        RECT 42.845 183.785 43.015 183.955 ;
        RECT 43.305 183.785 43.475 183.955 ;
        RECT 43.765 183.785 43.935 183.955 ;
        RECT 44.225 183.785 44.395 183.955 ;
        RECT 44.685 183.785 44.855 183.955 ;
        RECT 45.145 183.785 45.315 183.955 ;
        RECT 45.605 183.785 45.775 183.955 ;
        RECT 46.065 183.785 46.235 183.955 ;
        RECT 46.525 183.785 46.695 183.955 ;
        RECT 46.985 183.785 47.155 183.955 ;
        RECT 47.445 183.785 47.615 183.955 ;
        RECT 47.905 183.785 48.075 183.955 ;
        RECT 48.365 183.785 48.535 183.955 ;
        RECT 48.825 183.785 48.995 183.955 ;
        RECT 49.285 183.785 49.455 183.955 ;
        RECT 49.745 183.785 49.915 183.955 ;
        RECT 50.205 183.785 50.375 183.955 ;
        RECT 50.665 183.785 50.835 183.955 ;
        RECT 51.125 183.785 51.295 183.955 ;
        RECT 51.585 183.785 51.755 183.955 ;
        RECT 52.045 183.785 52.215 183.955 ;
        RECT 52.505 183.785 52.675 183.955 ;
        RECT 52.965 183.785 53.135 183.955 ;
        RECT 53.425 183.785 53.595 183.955 ;
        RECT 53.885 183.785 54.055 183.955 ;
        RECT 54.345 183.785 54.515 183.955 ;
        RECT 54.805 183.785 54.975 183.955 ;
        RECT 55.265 183.785 55.435 183.955 ;
        RECT 55.725 183.785 55.895 183.955 ;
        RECT 56.185 183.785 56.355 183.955 ;
        RECT 56.645 183.785 56.815 183.955 ;
        RECT 57.105 183.785 57.275 183.955 ;
        RECT 57.565 183.785 57.735 183.955 ;
        RECT 58.025 183.785 58.195 183.955 ;
        RECT 58.485 183.785 58.655 183.955 ;
        RECT 58.945 183.785 59.115 183.955 ;
        RECT 59.405 183.785 59.575 183.955 ;
        RECT 59.865 183.785 60.035 183.955 ;
        RECT 60.325 183.785 60.495 183.955 ;
        RECT 60.785 183.785 60.955 183.955 ;
        RECT 61.245 183.785 61.415 183.955 ;
        RECT 61.705 183.785 61.875 183.955 ;
        RECT 62.165 183.785 62.335 183.955 ;
        RECT 62.625 183.785 62.795 183.955 ;
        RECT 63.085 183.785 63.255 183.955 ;
        RECT 63.545 183.785 63.715 183.955 ;
        RECT 64.005 183.785 64.175 183.955 ;
        RECT 64.465 183.785 64.635 183.955 ;
        RECT 64.925 183.785 65.095 183.955 ;
        RECT 65.385 183.785 65.555 183.955 ;
        RECT 65.845 183.785 66.015 183.955 ;
        RECT 66.305 183.785 66.475 183.955 ;
        RECT 66.765 183.785 66.935 183.955 ;
        RECT 67.225 183.785 67.395 183.955 ;
        RECT 67.685 183.785 67.855 183.955 ;
        RECT 68.145 183.785 68.315 183.955 ;
        RECT 68.605 183.785 68.775 183.955 ;
        RECT 69.065 183.785 69.235 183.955 ;
        RECT 69.525 183.785 69.695 183.955 ;
        RECT 69.985 183.785 70.155 183.955 ;
        RECT 70.445 183.785 70.615 183.955 ;
        RECT 70.905 183.785 71.075 183.955 ;
        RECT 71.365 183.785 71.535 183.955 ;
        RECT 71.825 183.785 71.995 183.955 ;
        RECT 72.285 183.785 72.455 183.955 ;
        RECT 72.745 183.785 72.915 183.955 ;
        RECT 73.205 183.785 73.375 183.955 ;
        RECT 73.665 183.785 73.835 183.955 ;
        RECT 74.125 183.785 74.295 183.955 ;
        RECT 74.585 183.785 74.755 183.955 ;
        RECT 75.045 183.785 75.215 183.955 ;
        RECT 75.505 183.785 75.675 183.955 ;
        RECT 75.965 183.785 76.135 183.955 ;
        RECT 76.425 183.785 76.595 183.955 ;
        RECT 76.885 183.785 77.055 183.955 ;
        RECT 77.345 183.785 77.515 183.955 ;
        RECT 77.805 183.785 77.975 183.955 ;
        RECT 78.265 183.785 78.435 183.955 ;
        RECT 78.725 183.785 78.895 183.955 ;
        RECT 79.185 183.785 79.355 183.955 ;
        RECT 79.645 183.785 79.815 183.955 ;
        RECT 80.105 183.785 80.275 183.955 ;
        RECT 80.565 183.785 80.735 183.955 ;
        RECT 81.025 183.785 81.195 183.955 ;
        RECT 81.485 183.785 81.655 183.955 ;
        RECT 81.945 183.785 82.115 183.955 ;
        RECT 82.405 183.785 82.575 183.955 ;
        RECT 82.865 183.785 83.035 183.955 ;
        RECT 83.325 183.785 83.495 183.955 ;
        RECT 83.785 183.785 83.955 183.955 ;
        RECT 84.245 183.785 84.415 183.955 ;
        RECT 84.705 183.785 84.875 183.955 ;
        RECT 85.165 183.785 85.335 183.955 ;
        RECT 85.625 183.785 85.795 183.955 ;
        RECT 86.085 183.785 86.255 183.955 ;
        RECT 86.545 183.785 86.715 183.955 ;
        RECT 87.005 183.785 87.175 183.955 ;
        RECT 87.465 183.785 87.635 183.955 ;
        RECT 87.925 183.785 88.095 183.955 ;
        RECT 88.385 183.785 88.555 183.955 ;
        RECT 88.845 183.785 89.015 183.955 ;
        RECT 89.305 183.785 89.475 183.955 ;
        RECT 89.765 183.785 89.935 183.955 ;
        RECT 90.225 183.785 90.395 183.955 ;
        RECT 90.685 183.785 90.855 183.955 ;
        RECT 91.145 183.785 91.315 183.955 ;
        RECT 91.605 183.785 91.775 183.955 ;
        RECT 92.065 183.785 92.235 183.955 ;
        RECT 92.525 183.785 92.695 183.955 ;
        RECT 92.985 183.785 93.155 183.955 ;
        RECT 93.445 183.785 93.615 183.955 ;
        RECT 93.905 183.785 94.075 183.955 ;
        RECT 94.365 183.785 94.535 183.955 ;
        RECT 94.825 183.785 94.995 183.955 ;
        RECT 95.285 183.785 95.455 183.955 ;
        RECT 95.745 183.785 95.915 183.955 ;
        RECT 96.205 183.785 96.375 183.955 ;
        RECT 96.665 183.785 96.835 183.955 ;
        RECT 97.125 183.785 97.295 183.955 ;
        RECT 97.585 183.785 97.755 183.955 ;
        RECT 98.045 183.785 98.215 183.955 ;
        RECT 98.505 183.785 98.675 183.955 ;
        RECT 98.965 183.785 99.135 183.955 ;
        RECT 99.425 183.785 99.595 183.955 ;
        RECT 99.885 183.785 100.055 183.955 ;
        RECT 100.345 183.785 100.515 183.955 ;
        RECT 100.805 183.785 100.975 183.955 ;
        RECT 101.265 183.785 101.435 183.955 ;
        RECT 101.725 183.785 101.895 183.955 ;
        RECT 102.185 183.785 102.355 183.955 ;
        RECT 102.645 183.785 102.815 183.955 ;
        RECT 103.105 183.785 103.275 183.955 ;
        RECT 103.565 183.785 103.735 183.955 ;
        RECT 104.025 183.785 104.195 183.955 ;
        RECT 104.485 183.785 104.655 183.955 ;
        RECT 104.945 183.785 105.115 183.955 ;
        RECT 105.405 183.785 105.575 183.955 ;
        RECT 105.865 183.785 106.035 183.955 ;
        RECT 106.325 183.785 106.495 183.955 ;
        RECT 106.785 183.785 106.955 183.955 ;
        RECT 107.245 183.785 107.415 183.955 ;
        RECT 107.705 183.785 107.875 183.955 ;
        RECT 108.165 183.785 108.335 183.955 ;
        RECT 108.625 183.785 108.795 183.955 ;
        RECT 109.085 183.785 109.255 183.955 ;
        RECT 109.545 183.785 109.715 183.955 ;
        RECT 110.005 183.785 110.175 183.955 ;
        RECT 110.465 183.785 110.635 183.955 ;
        RECT 110.925 183.785 111.095 183.955 ;
        RECT 111.385 183.785 111.555 183.955 ;
        RECT 111.845 183.785 112.015 183.955 ;
        RECT 112.305 183.785 112.475 183.955 ;
        RECT 112.765 183.785 112.935 183.955 ;
        RECT 113.225 183.785 113.395 183.955 ;
        RECT 113.685 183.785 113.855 183.955 ;
        RECT 114.145 183.785 114.315 183.955 ;
        RECT 114.605 183.785 114.775 183.955 ;
        RECT 115.065 183.785 115.235 183.955 ;
        RECT 115.525 183.785 115.695 183.955 ;
        RECT 41.925 178.345 42.095 178.515 ;
        RECT 42.385 178.345 42.555 178.515 ;
        RECT 42.845 178.345 43.015 178.515 ;
        RECT 43.305 178.345 43.475 178.515 ;
        RECT 43.765 178.345 43.935 178.515 ;
        RECT 44.225 178.345 44.395 178.515 ;
        RECT 44.685 178.345 44.855 178.515 ;
        RECT 45.145 178.345 45.315 178.515 ;
        RECT 45.605 178.345 45.775 178.515 ;
        RECT 46.065 178.345 46.235 178.515 ;
        RECT 46.525 178.345 46.695 178.515 ;
        RECT 46.985 178.345 47.155 178.515 ;
        RECT 47.445 178.345 47.615 178.515 ;
        RECT 47.905 178.345 48.075 178.515 ;
        RECT 48.365 178.345 48.535 178.515 ;
        RECT 48.825 178.345 48.995 178.515 ;
        RECT 49.285 178.345 49.455 178.515 ;
        RECT 49.745 178.345 49.915 178.515 ;
        RECT 50.205 178.345 50.375 178.515 ;
        RECT 50.665 178.345 50.835 178.515 ;
        RECT 51.125 178.345 51.295 178.515 ;
        RECT 51.585 178.345 51.755 178.515 ;
        RECT 52.045 178.345 52.215 178.515 ;
        RECT 52.505 178.345 52.675 178.515 ;
        RECT 52.965 178.345 53.135 178.515 ;
        RECT 53.425 178.345 53.595 178.515 ;
        RECT 53.885 178.345 54.055 178.515 ;
        RECT 54.345 178.345 54.515 178.515 ;
        RECT 54.805 178.345 54.975 178.515 ;
        RECT 55.265 178.345 55.435 178.515 ;
        RECT 55.725 178.345 55.895 178.515 ;
        RECT 56.185 178.345 56.355 178.515 ;
        RECT 56.645 178.345 56.815 178.515 ;
        RECT 57.105 178.345 57.275 178.515 ;
        RECT 57.565 178.345 57.735 178.515 ;
        RECT 58.025 178.345 58.195 178.515 ;
        RECT 58.485 178.345 58.655 178.515 ;
        RECT 58.945 178.345 59.115 178.515 ;
        RECT 59.405 178.345 59.575 178.515 ;
        RECT 59.865 178.345 60.035 178.515 ;
        RECT 60.325 178.345 60.495 178.515 ;
        RECT 60.785 178.345 60.955 178.515 ;
        RECT 61.245 178.345 61.415 178.515 ;
        RECT 61.705 178.345 61.875 178.515 ;
        RECT 62.165 178.345 62.335 178.515 ;
        RECT 62.625 178.345 62.795 178.515 ;
        RECT 63.085 178.345 63.255 178.515 ;
        RECT 63.545 178.345 63.715 178.515 ;
        RECT 64.005 178.345 64.175 178.515 ;
        RECT 64.465 178.345 64.635 178.515 ;
        RECT 64.925 178.345 65.095 178.515 ;
        RECT 65.385 178.345 65.555 178.515 ;
        RECT 65.845 178.345 66.015 178.515 ;
        RECT 66.305 178.345 66.475 178.515 ;
        RECT 66.765 178.345 66.935 178.515 ;
        RECT 67.225 178.345 67.395 178.515 ;
        RECT 67.685 178.345 67.855 178.515 ;
        RECT 68.145 178.345 68.315 178.515 ;
        RECT 68.605 178.345 68.775 178.515 ;
        RECT 69.065 178.345 69.235 178.515 ;
        RECT 69.525 178.345 69.695 178.515 ;
        RECT 69.985 178.345 70.155 178.515 ;
        RECT 70.445 178.345 70.615 178.515 ;
        RECT 70.905 178.345 71.075 178.515 ;
        RECT 71.365 178.345 71.535 178.515 ;
        RECT 71.825 178.345 71.995 178.515 ;
        RECT 72.285 178.345 72.455 178.515 ;
        RECT 72.745 178.345 72.915 178.515 ;
        RECT 73.205 178.345 73.375 178.515 ;
        RECT 73.665 178.345 73.835 178.515 ;
        RECT 74.125 178.345 74.295 178.515 ;
        RECT 74.585 178.345 74.755 178.515 ;
        RECT 75.045 178.345 75.215 178.515 ;
        RECT 75.505 178.345 75.675 178.515 ;
        RECT 75.965 178.345 76.135 178.515 ;
        RECT 76.425 178.345 76.595 178.515 ;
        RECT 76.885 178.345 77.055 178.515 ;
        RECT 77.345 178.345 77.515 178.515 ;
        RECT 77.805 178.345 77.975 178.515 ;
        RECT 78.265 178.345 78.435 178.515 ;
        RECT 78.725 178.345 78.895 178.515 ;
        RECT 79.185 178.345 79.355 178.515 ;
        RECT 79.645 178.345 79.815 178.515 ;
        RECT 80.105 178.345 80.275 178.515 ;
        RECT 80.565 178.345 80.735 178.515 ;
        RECT 81.025 178.345 81.195 178.515 ;
        RECT 81.485 178.345 81.655 178.515 ;
        RECT 81.945 178.345 82.115 178.515 ;
        RECT 82.405 178.345 82.575 178.515 ;
        RECT 82.865 178.345 83.035 178.515 ;
        RECT 83.325 178.345 83.495 178.515 ;
        RECT 83.785 178.345 83.955 178.515 ;
        RECT 84.245 178.345 84.415 178.515 ;
        RECT 84.705 178.345 84.875 178.515 ;
        RECT 85.165 178.345 85.335 178.515 ;
        RECT 85.625 178.345 85.795 178.515 ;
        RECT 86.085 178.345 86.255 178.515 ;
        RECT 86.545 178.345 86.715 178.515 ;
        RECT 87.005 178.345 87.175 178.515 ;
        RECT 87.465 178.345 87.635 178.515 ;
        RECT 87.925 178.345 88.095 178.515 ;
        RECT 88.385 178.345 88.555 178.515 ;
        RECT 88.845 178.345 89.015 178.515 ;
        RECT 89.305 178.345 89.475 178.515 ;
        RECT 89.765 178.345 89.935 178.515 ;
        RECT 90.225 178.345 90.395 178.515 ;
        RECT 90.685 178.345 90.855 178.515 ;
        RECT 91.145 178.345 91.315 178.515 ;
        RECT 91.605 178.345 91.775 178.515 ;
        RECT 92.065 178.345 92.235 178.515 ;
        RECT 92.525 178.345 92.695 178.515 ;
        RECT 92.985 178.345 93.155 178.515 ;
        RECT 93.445 178.345 93.615 178.515 ;
        RECT 93.905 178.345 94.075 178.515 ;
        RECT 94.365 178.345 94.535 178.515 ;
        RECT 94.825 178.345 94.995 178.515 ;
        RECT 95.285 178.345 95.455 178.515 ;
        RECT 95.745 178.345 95.915 178.515 ;
        RECT 96.205 178.345 96.375 178.515 ;
        RECT 96.665 178.345 96.835 178.515 ;
        RECT 97.125 178.345 97.295 178.515 ;
        RECT 97.585 178.345 97.755 178.515 ;
        RECT 98.045 178.345 98.215 178.515 ;
        RECT 98.505 178.345 98.675 178.515 ;
        RECT 98.965 178.345 99.135 178.515 ;
        RECT 99.425 178.345 99.595 178.515 ;
        RECT 99.885 178.345 100.055 178.515 ;
        RECT 100.345 178.345 100.515 178.515 ;
        RECT 100.805 178.345 100.975 178.515 ;
        RECT 101.265 178.345 101.435 178.515 ;
        RECT 101.725 178.345 101.895 178.515 ;
        RECT 102.185 178.345 102.355 178.515 ;
        RECT 102.645 178.345 102.815 178.515 ;
        RECT 103.105 178.345 103.275 178.515 ;
        RECT 103.565 178.345 103.735 178.515 ;
        RECT 104.025 178.345 104.195 178.515 ;
        RECT 104.485 178.345 104.655 178.515 ;
        RECT 104.945 178.345 105.115 178.515 ;
        RECT 105.405 178.345 105.575 178.515 ;
        RECT 105.865 178.345 106.035 178.515 ;
        RECT 106.325 178.345 106.495 178.515 ;
        RECT 106.785 178.345 106.955 178.515 ;
        RECT 107.245 178.345 107.415 178.515 ;
        RECT 107.705 178.345 107.875 178.515 ;
        RECT 108.165 178.345 108.335 178.515 ;
        RECT 108.625 178.345 108.795 178.515 ;
        RECT 109.085 178.345 109.255 178.515 ;
        RECT 109.545 178.345 109.715 178.515 ;
        RECT 110.005 178.345 110.175 178.515 ;
        RECT 110.465 178.345 110.635 178.515 ;
        RECT 110.925 178.345 111.095 178.515 ;
        RECT 111.385 178.345 111.555 178.515 ;
        RECT 111.845 178.345 112.015 178.515 ;
        RECT 112.305 178.345 112.475 178.515 ;
        RECT 112.765 178.345 112.935 178.515 ;
        RECT 113.225 178.345 113.395 178.515 ;
        RECT 113.685 178.345 113.855 178.515 ;
        RECT 114.145 178.345 114.315 178.515 ;
        RECT 114.605 178.345 114.775 178.515 ;
        RECT 115.065 178.345 115.235 178.515 ;
        RECT 115.525 178.345 115.695 178.515 ;
        RECT 41.925 172.905 42.095 173.075 ;
        RECT 42.385 172.905 42.555 173.075 ;
        RECT 42.845 172.905 43.015 173.075 ;
        RECT 43.305 172.905 43.475 173.075 ;
        RECT 43.765 172.905 43.935 173.075 ;
        RECT 44.225 172.905 44.395 173.075 ;
        RECT 44.685 172.905 44.855 173.075 ;
        RECT 45.145 172.905 45.315 173.075 ;
        RECT 45.605 172.905 45.775 173.075 ;
        RECT 46.065 172.905 46.235 173.075 ;
        RECT 46.525 172.905 46.695 173.075 ;
        RECT 46.985 172.905 47.155 173.075 ;
        RECT 47.445 172.905 47.615 173.075 ;
        RECT 47.905 172.905 48.075 173.075 ;
        RECT 48.365 172.905 48.535 173.075 ;
        RECT 48.825 172.905 48.995 173.075 ;
        RECT 49.285 172.905 49.455 173.075 ;
        RECT 49.745 172.905 49.915 173.075 ;
        RECT 50.205 172.905 50.375 173.075 ;
        RECT 50.665 172.905 50.835 173.075 ;
        RECT 51.125 172.905 51.295 173.075 ;
        RECT 51.585 172.905 51.755 173.075 ;
        RECT 52.045 172.905 52.215 173.075 ;
        RECT 52.505 172.905 52.675 173.075 ;
        RECT 52.965 172.905 53.135 173.075 ;
        RECT 53.425 172.905 53.595 173.075 ;
        RECT 53.885 172.905 54.055 173.075 ;
        RECT 54.345 172.905 54.515 173.075 ;
        RECT 54.805 172.905 54.975 173.075 ;
        RECT 55.265 172.905 55.435 173.075 ;
        RECT 55.725 172.905 55.895 173.075 ;
        RECT 56.185 172.905 56.355 173.075 ;
        RECT 56.645 172.905 56.815 173.075 ;
        RECT 57.105 172.905 57.275 173.075 ;
        RECT 57.565 172.905 57.735 173.075 ;
        RECT 58.025 172.905 58.195 173.075 ;
        RECT 58.485 172.905 58.655 173.075 ;
        RECT 58.945 172.905 59.115 173.075 ;
        RECT 59.405 172.905 59.575 173.075 ;
        RECT 59.865 172.905 60.035 173.075 ;
        RECT 60.325 172.905 60.495 173.075 ;
        RECT 60.785 172.905 60.955 173.075 ;
        RECT 61.245 172.905 61.415 173.075 ;
        RECT 61.705 172.905 61.875 173.075 ;
        RECT 62.165 172.905 62.335 173.075 ;
        RECT 62.625 172.905 62.795 173.075 ;
        RECT 63.085 172.905 63.255 173.075 ;
        RECT 63.545 172.905 63.715 173.075 ;
        RECT 64.005 172.905 64.175 173.075 ;
        RECT 64.465 172.905 64.635 173.075 ;
        RECT 64.925 172.905 65.095 173.075 ;
        RECT 65.385 172.905 65.555 173.075 ;
        RECT 65.845 172.905 66.015 173.075 ;
        RECT 66.305 172.905 66.475 173.075 ;
        RECT 66.765 172.905 66.935 173.075 ;
        RECT 67.225 172.905 67.395 173.075 ;
        RECT 67.685 172.905 67.855 173.075 ;
        RECT 68.145 172.905 68.315 173.075 ;
        RECT 68.605 172.905 68.775 173.075 ;
        RECT 69.065 172.905 69.235 173.075 ;
        RECT 69.525 172.905 69.695 173.075 ;
        RECT 69.985 172.905 70.155 173.075 ;
        RECT 70.445 172.905 70.615 173.075 ;
        RECT 70.905 172.905 71.075 173.075 ;
        RECT 71.365 172.905 71.535 173.075 ;
        RECT 71.825 172.905 71.995 173.075 ;
        RECT 72.285 172.905 72.455 173.075 ;
        RECT 72.745 172.905 72.915 173.075 ;
        RECT 73.205 172.905 73.375 173.075 ;
        RECT 73.665 172.905 73.835 173.075 ;
        RECT 74.125 172.905 74.295 173.075 ;
        RECT 74.585 172.905 74.755 173.075 ;
        RECT 75.045 172.905 75.215 173.075 ;
        RECT 75.505 172.905 75.675 173.075 ;
        RECT 75.965 172.905 76.135 173.075 ;
        RECT 76.425 172.905 76.595 173.075 ;
        RECT 76.885 172.905 77.055 173.075 ;
        RECT 77.345 172.905 77.515 173.075 ;
        RECT 77.805 172.905 77.975 173.075 ;
        RECT 78.265 172.905 78.435 173.075 ;
        RECT 78.725 172.905 78.895 173.075 ;
        RECT 79.185 172.905 79.355 173.075 ;
        RECT 79.645 172.905 79.815 173.075 ;
        RECT 80.105 172.905 80.275 173.075 ;
        RECT 80.565 172.905 80.735 173.075 ;
        RECT 81.025 172.905 81.195 173.075 ;
        RECT 81.485 172.905 81.655 173.075 ;
        RECT 81.945 172.905 82.115 173.075 ;
        RECT 82.405 172.905 82.575 173.075 ;
        RECT 82.865 172.905 83.035 173.075 ;
        RECT 83.325 172.905 83.495 173.075 ;
        RECT 83.785 172.905 83.955 173.075 ;
        RECT 84.245 172.905 84.415 173.075 ;
        RECT 84.705 172.905 84.875 173.075 ;
        RECT 85.165 172.905 85.335 173.075 ;
        RECT 85.625 172.905 85.795 173.075 ;
        RECT 86.085 172.905 86.255 173.075 ;
        RECT 86.545 172.905 86.715 173.075 ;
        RECT 87.005 172.905 87.175 173.075 ;
        RECT 87.465 172.905 87.635 173.075 ;
        RECT 87.925 172.905 88.095 173.075 ;
        RECT 88.385 172.905 88.555 173.075 ;
        RECT 88.845 172.905 89.015 173.075 ;
        RECT 89.305 172.905 89.475 173.075 ;
        RECT 89.765 172.905 89.935 173.075 ;
        RECT 90.225 172.905 90.395 173.075 ;
        RECT 90.685 172.905 90.855 173.075 ;
        RECT 91.145 172.905 91.315 173.075 ;
        RECT 91.605 172.905 91.775 173.075 ;
        RECT 92.065 172.905 92.235 173.075 ;
        RECT 92.525 172.905 92.695 173.075 ;
        RECT 92.985 172.905 93.155 173.075 ;
        RECT 93.445 172.905 93.615 173.075 ;
        RECT 93.905 172.905 94.075 173.075 ;
        RECT 94.365 172.905 94.535 173.075 ;
        RECT 94.825 172.905 94.995 173.075 ;
        RECT 95.285 172.905 95.455 173.075 ;
        RECT 95.745 172.905 95.915 173.075 ;
        RECT 96.205 172.905 96.375 173.075 ;
        RECT 96.665 172.905 96.835 173.075 ;
        RECT 97.125 172.905 97.295 173.075 ;
        RECT 97.585 172.905 97.755 173.075 ;
        RECT 98.045 172.905 98.215 173.075 ;
        RECT 98.505 172.905 98.675 173.075 ;
        RECT 98.965 172.905 99.135 173.075 ;
        RECT 99.425 172.905 99.595 173.075 ;
        RECT 99.885 172.905 100.055 173.075 ;
        RECT 100.345 172.905 100.515 173.075 ;
        RECT 100.805 172.905 100.975 173.075 ;
        RECT 101.265 172.905 101.435 173.075 ;
        RECT 101.725 172.905 101.895 173.075 ;
        RECT 102.185 172.905 102.355 173.075 ;
        RECT 102.645 172.905 102.815 173.075 ;
        RECT 103.105 172.905 103.275 173.075 ;
        RECT 103.565 172.905 103.735 173.075 ;
        RECT 104.025 172.905 104.195 173.075 ;
        RECT 104.485 172.905 104.655 173.075 ;
        RECT 104.945 172.905 105.115 173.075 ;
        RECT 105.405 172.905 105.575 173.075 ;
        RECT 105.865 172.905 106.035 173.075 ;
        RECT 106.325 172.905 106.495 173.075 ;
        RECT 106.785 172.905 106.955 173.075 ;
        RECT 107.245 172.905 107.415 173.075 ;
        RECT 107.705 172.905 107.875 173.075 ;
        RECT 108.165 172.905 108.335 173.075 ;
        RECT 108.625 172.905 108.795 173.075 ;
        RECT 109.085 172.905 109.255 173.075 ;
        RECT 109.545 172.905 109.715 173.075 ;
        RECT 110.005 172.905 110.175 173.075 ;
        RECT 110.465 172.905 110.635 173.075 ;
        RECT 110.925 172.905 111.095 173.075 ;
        RECT 111.385 172.905 111.555 173.075 ;
        RECT 111.845 172.905 112.015 173.075 ;
        RECT 112.305 172.905 112.475 173.075 ;
        RECT 112.765 172.905 112.935 173.075 ;
        RECT 113.225 172.905 113.395 173.075 ;
        RECT 113.685 172.905 113.855 173.075 ;
        RECT 114.145 172.905 114.315 173.075 ;
        RECT 114.605 172.905 114.775 173.075 ;
        RECT 115.065 172.905 115.235 173.075 ;
        RECT 115.525 172.905 115.695 173.075 ;
        RECT 41.925 167.465 42.095 167.635 ;
        RECT 42.385 167.465 42.555 167.635 ;
        RECT 42.845 167.465 43.015 167.635 ;
        RECT 43.305 167.465 43.475 167.635 ;
        RECT 43.765 167.465 43.935 167.635 ;
        RECT 44.225 167.465 44.395 167.635 ;
        RECT 44.685 167.465 44.855 167.635 ;
        RECT 45.145 167.465 45.315 167.635 ;
        RECT 45.605 167.465 45.775 167.635 ;
        RECT 46.065 167.465 46.235 167.635 ;
        RECT 46.525 167.465 46.695 167.635 ;
        RECT 46.985 167.465 47.155 167.635 ;
        RECT 47.445 167.465 47.615 167.635 ;
        RECT 47.905 167.465 48.075 167.635 ;
        RECT 48.365 167.465 48.535 167.635 ;
        RECT 48.825 167.465 48.995 167.635 ;
        RECT 49.285 167.465 49.455 167.635 ;
        RECT 49.745 167.465 49.915 167.635 ;
        RECT 50.205 167.465 50.375 167.635 ;
        RECT 50.665 167.465 50.835 167.635 ;
        RECT 51.125 167.465 51.295 167.635 ;
        RECT 51.585 167.465 51.755 167.635 ;
        RECT 52.045 167.465 52.215 167.635 ;
        RECT 52.505 167.465 52.675 167.635 ;
        RECT 52.965 167.465 53.135 167.635 ;
        RECT 53.425 167.465 53.595 167.635 ;
        RECT 53.885 167.465 54.055 167.635 ;
        RECT 54.345 167.465 54.515 167.635 ;
        RECT 54.805 167.465 54.975 167.635 ;
        RECT 55.265 167.465 55.435 167.635 ;
        RECT 55.725 167.465 55.895 167.635 ;
        RECT 56.185 167.465 56.355 167.635 ;
        RECT 56.645 167.465 56.815 167.635 ;
        RECT 57.105 167.465 57.275 167.635 ;
        RECT 57.565 167.465 57.735 167.635 ;
        RECT 58.025 167.465 58.195 167.635 ;
        RECT 58.485 167.465 58.655 167.635 ;
        RECT 58.945 167.465 59.115 167.635 ;
        RECT 59.405 167.465 59.575 167.635 ;
        RECT 59.865 167.465 60.035 167.635 ;
        RECT 60.325 167.465 60.495 167.635 ;
        RECT 60.785 167.465 60.955 167.635 ;
        RECT 61.245 167.465 61.415 167.635 ;
        RECT 61.705 167.465 61.875 167.635 ;
        RECT 62.165 167.465 62.335 167.635 ;
        RECT 62.625 167.465 62.795 167.635 ;
        RECT 63.085 167.465 63.255 167.635 ;
        RECT 63.545 167.465 63.715 167.635 ;
        RECT 64.005 167.465 64.175 167.635 ;
        RECT 64.465 167.465 64.635 167.635 ;
        RECT 64.925 167.465 65.095 167.635 ;
        RECT 65.385 167.465 65.555 167.635 ;
        RECT 65.845 167.465 66.015 167.635 ;
        RECT 66.305 167.465 66.475 167.635 ;
        RECT 66.765 167.465 66.935 167.635 ;
        RECT 67.225 167.465 67.395 167.635 ;
        RECT 67.685 167.465 67.855 167.635 ;
        RECT 68.145 167.465 68.315 167.635 ;
        RECT 68.605 167.465 68.775 167.635 ;
        RECT 69.065 167.465 69.235 167.635 ;
        RECT 69.525 167.465 69.695 167.635 ;
        RECT 69.985 167.465 70.155 167.635 ;
        RECT 70.445 167.465 70.615 167.635 ;
        RECT 70.905 167.465 71.075 167.635 ;
        RECT 71.365 167.465 71.535 167.635 ;
        RECT 71.825 167.465 71.995 167.635 ;
        RECT 72.285 167.465 72.455 167.635 ;
        RECT 72.745 167.465 72.915 167.635 ;
        RECT 73.205 167.465 73.375 167.635 ;
        RECT 73.665 167.465 73.835 167.635 ;
        RECT 74.125 167.465 74.295 167.635 ;
        RECT 74.585 167.465 74.755 167.635 ;
        RECT 75.045 167.465 75.215 167.635 ;
        RECT 75.505 167.465 75.675 167.635 ;
        RECT 75.965 167.465 76.135 167.635 ;
        RECT 76.425 167.465 76.595 167.635 ;
        RECT 76.885 167.465 77.055 167.635 ;
        RECT 77.345 167.465 77.515 167.635 ;
        RECT 77.805 167.465 77.975 167.635 ;
        RECT 78.265 167.465 78.435 167.635 ;
        RECT 78.725 167.465 78.895 167.635 ;
        RECT 79.185 167.465 79.355 167.635 ;
        RECT 79.645 167.465 79.815 167.635 ;
        RECT 80.105 167.465 80.275 167.635 ;
        RECT 80.565 167.465 80.735 167.635 ;
        RECT 81.025 167.465 81.195 167.635 ;
        RECT 81.485 167.465 81.655 167.635 ;
        RECT 81.945 167.465 82.115 167.635 ;
        RECT 82.405 167.465 82.575 167.635 ;
        RECT 82.865 167.465 83.035 167.635 ;
        RECT 83.325 167.465 83.495 167.635 ;
        RECT 83.785 167.465 83.955 167.635 ;
        RECT 84.245 167.465 84.415 167.635 ;
        RECT 84.705 167.465 84.875 167.635 ;
        RECT 85.165 167.465 85.335 167.635 ;
        RECT 85.625 167.465 85.795 167.635 ;
        RECT 86.085 167.465 86.255 167.635 ;
        RECT 86.545 167.465 86.715 167.635 ;
        RECT 87.005 167.465 87.175 167.635 ;
        RECT 87.465 167.465 87.635 167.635 ;
        RECT 87.925 167.465 88.095 167.635 ;
        RECT 88.385 167.465 88.555 167.635 ;
        RECT 88.845 167.465 89.015 167.635 ;
        RECT 89.305 167.465 89.475 167.635 ;
        RECT 89.765 167.465 89.935 167.635 ;
        RECT 90.225 167.465 90.395 167.635 ;
        RECT 90.685 167.465 90.855 167.635 ;
        RECT 91.145 167.465 91.315 167.635 ;
        RECT 91.605 167.465 91.775 167.635 ;
        RECT 92.065 167.465 92.235 167.635 ;
        RECT 92.525 167.465 92.695 167.635 ;
        RECT 92.985 167.465 93.155 167.635 ;
        RECT 93.445 167.465 93.615 167.635 ;
        RECT 93.905 167.465 94.075 167.635 ;
        RECT 94.365 167.465 94.535 167.635 ;
        RECT 94.825 167.465 94.995 167.635 ;
        RECT 95.285 167.465 95.455 167.635 ;
        RECT 95.745 167.465 95.915 167.635 ;
        RECT 96.205 167.465 96.375 167.635 ;
        RECT 96.665 167.465 96.835 167.635 ;
        RECT 97.125 167.465 97.295 167.635 ;
        RECT 97.585 167.465 97.755 167.635 ;
        RECT 98.045 167.465 98.215 167.635 ;
        RECT 98.505 167.465 98.675 167.635 ;
        RECT 98.965 167.465 99.135 167.635 ;
        RECT 99.425 167.465 99.595 167.635 ;
        RECT 99.885 167.465 100.055 167.635 ;
        RECT 100.345 167.465 100.515 167.635 ;
        RECT 100.805 167.465 100.975 167.635 ;
        RECT 101.265 167.465 101.435 167.635 ;
        RECT 101.725 167.465 101.895 167.635 ;
        RECT 102.185 167.465 102.355 167.635 ;
        RECT 102.645 167.465 102.815 167.635 ;
        RECT 103.105 167.465 103.275 167.635 ;
        RECT 103.565 167.465 103.735 167.635 ;
        RECT 104.025 167.465 104.195 167.635 ;
        RECT 104.485 167.465 104.655 167.635 ;
        RECT 104.945 167.465 105.115 167.635 ;
        RECT 105.405 167.465 105.575 167.635 ;
        RECT 105.865 167.465 106.035 167.635 ;
        RECT 106.325 167.465 106.495 167.635 ;
        RECT 106.785 167.465 106.955 167.635 ;
        RECT 107.245 167.465 107.415 167.635 ;
        RECT 107.705 167.465 107.875 167.635 ;
        RECT 108.165 167.465 108.335 167.635 ;
        RECT 108.625 167.465 108.795 167.635 ;
        RECT 109.085 167.465 109.255 167.635 ;
        RECT 109.545 167.465 109.715 167.635 ;
        RECT 110.005 167.465 110.175 167.635 ;
        RECT 110.465 167.465 110.635 167.635 ;
        RECT 110.925 167.465 111.095 167.635 ;
        RECT 111.385 167.465 111.555 167.635 ;
        RECT 111.845 167.465 112.015 167.635 ;
        RECT 112.305 167.465 112.475 167.635 ;
        RECT 112.765 167.465 112.935 167.635 ;
        RECT 113.225 167.465 113.395 167.635 ;
        RECT 113.685 167.465 113.855 167.635 ;
        RECT 114.145 167.465 114.315 167.635 ;
        RECT 114.605 167.465 114.775 167.635 ;
        RECT 115.065 167.465 115.235 167.635 ;
        RECT 115.525 167.465 115.695 167.635 ;
        RECT 41.925 162.025 42.095 162.195 ;
        RECT 42.385 162.025 42.555 162.195 ;
        RECT 42.845 162.025 43.015 162.195 ;
        RECT 43.305 162.025 43.475 162.195 ;
        RECT 43.765 162.025 43.935 162.195 ;
        RECT 44.225 162.025 44.395 162.195 ;
        RECT 44.685 162.025 44.855 162.195 ;
        RECT 45.145 162.025 45.315 162.195 ;
        RECT 45.605 162.025 45.775 162.195 ;
        RECT 46.065 162.025 46.235 162.195 ;
        RECT 46.525 162.025 46.695 162.195 ;
        RECT 46.985 162.025 47.155 162.195 ;
        RECT 47.445 162.025 47.615 162.195 ;
        RECT 47.905 162.025 48.075 162.195 ;
        RECT 48.365 162.025 48.535 162.195 ;
        RECT 48.825 162.025 48.995 162.195 ;
        RECT 49.285 162.025 49.455 162.195 ;
        RECT 49.745 162.025 49.915 162.195 ;
        RECT 50.205 162.025 50.375 162.195 ;
        RECT 50.665 162.025 50.835 162.195 ;
        RECT 51.125 162.025 51.295 162.195 ;
        RECT 51.585 162.025 51.755 162.195 ;
        RECT 52.045 162.025 52.215 162.195 ;
        RECT 52.505 162.025 52.675 162.195 ;
        RECT 52.965 162.025 53.135 162.195 ;
        RECT 53.425 162.025 53.595 162.195 ;
        RECT 53.885 162.025 54.055 162.195 ;
        RECT 54.345 162.025 54.515 162.195 ;
        RECT 54.805 162.025 54.975 162.195 ;
        RECT 55.265 162.025 55.435 162.195 ;
        RECT 55.725 162.025 55.895 162.195 ;
        RECT 56.185 162.025 56.355 162.195 ;
        RECT 56.645 162.025 56.815 162.195 ;
        RECT 57.105 162.025 57.275 162.195 ;
        RECT 57.565 162.025 57.735 162.195 ;
        RECT 58.025 162.025 58.195 162.195 ;
        RECT 58.485 162.025 58.655 162.195 ;
        RECT 58.945 162.025 59.115 162.195 ;
        RECT 59.405 162.025 59.575 162.195 ;
        RECT 59.865 162.025 60.035 162.195 ;
        RECT 60.325 162.025 60.495 162.195 ;
        RECT 60.785 162.025 60.955 162.195 ;
        RECT 61.245 162.025 61.415 162.195 ;
        RECT 61.705 162.025 61.875 162.195 ;
        RECT 62.165 162.025 62.335 162.195 ;
        RECT 62.625 162.025 62.795 162.195 ;
        RECT 63.085 162.025 63.255 162.195 ;
        RECT 63.545 162.025 63.715 162.195 ;
        RECT 64.005 162.025 64.175 162.195 ;
        RECT 64.465 162.025 64.635 162.195 ;
        RECT 64.925 162.025 65.095 162.195 ;
        RECT 65.385 162.025 65.555 162.195 ;
        RECT 65.845 162.025 66.015 162.195 ;
        RECT 66.305 162.025 66.475 162.195 ;
        RECT 66.765 162.025 66.935 162.195 ;
        RECT 67.225 162.025 67.395 162.195 ;
        RECT 67.685 162.025 67.855 162.195 ;
        RECT 68.145 162.025 68.315 162.195 ;
        RECT 68.605 162.025 68.775 162.195 ;
        RECT 69.065 162.025 69.235 162.195 ;
        RECT 69.525 162.025 69.695 162.195 ;
        RECT 69.985 162.025 70.155 162.195 ;
        RECT 70.445 162.025 70.615 162.195 ;
        RECT 70.905 162.025 71.075 162.195 ;
        RECT 71.365 162.025 71.535 162.195 ;
        RECT 71.825 162.025 71.995 162.195 ;
        RECT 72.285 162.025 72.455 162.195 ;
        RECT 72.745 162.025 72.915 162.195 ;
        RECT 73.205 162.025 73.375 162.195 ;
        RECT 73.665 162.025 73.835 162.195 ;
        RECT 74.125 162.025 74.295 162.195 ;
        RECT 74.585 162.025 74.755 162.195 ;
        RECT 75.045 162.025 75.215 162.195 ;
        RECT 75.505 162.025 75.675 162.195 ;
        RECT 75.965 162.025 76.135 162.195 ;
        RECT 76.425 162.025 76.595 162.195 ;
        RECT 76.885 162.025 77.055 162.195 ;
        RECT 77.345 162.025 77.515 162.195 ;
        RECT 77.805 162.025 77.975 162.195 ;
        RECT 78.265 162.025 78.435 162.195 ;
        RECT 78.725 162.025 78.895 162.195 ;
        RECT 79.185 162.025 79.355 162.195 ;
        RECT 79.645 162.025 79.815 162.195 ;
        RECT 80.105 162.025 80.275 162.195 ;
        RECT 80.565 162.025 80.735 162.195 ;
        RECT 81.025 162.025 81.195 162.195 ;
        RECT 81.485 162.025 81.655 162.195 ;
        RECT 81.945 162.025 82.115 162.195 ;
        RECT 82.405 162.025 82.575 162.195 ;
        RECT 82.865 162.025 83.035 162.195 ;
        RECT 83.325 162.025 83.495 162.195 ;
        RECT 83.785 162.025 83.955 162.195 ;
        RECT 84.245 162.025 84.415 162.195 ;
        RECT 84.705 162.025 84.875 162.195 ;
        RECT 85.165 162.025 85.335 162.195 ;
        RECT 85.625 162.025 85.795 162.195 ;
        RECT 86.085 162.025 86.255 162.195 ;
        RECT 86.545 162.025 86.715 162.195 ;
        RECT 87.005 162.025 87.175 162.195 ;
        RECT 87.465 162.025 87.635 162.195 ;
        RECT 87.925 162.025 88.095 162.195 ;
        RECT 88.385 162.025 88.555 162.195 ;
        RECT 88.845 162.025 89.015 162.195 ;
        RECT 89.305 162.025 89.475 162.195 ;
        RECT 89.765 162.025 89.935 162.195 ;
        RECT 90.225 162.025 90.395 162.195 ;
        RECT 90.685 162.025 90.855 162.195 ;
        RECT 91.145 162.025 91.315 162.195 ;
        RECT 91.605 162.025 91.775 162.195 ;
        RECT 92.065 162.025 92.235 162.195 ;
        RECT 92.525 162.025 92.695 162.195 ;
        RECT 92.985 162.025 93.155 162.195 ;
        RECT 93.445 162.025 93.615 162.195 ;
        RECT 93.905 162.025 94.075 162.195 ;
        RECT 94.365 162.025 94.535 162.195 ;
        RECT 94.825 162.025 94.995 162.195 ;
        RECT 95.285 162.025 95.455 162.195 ;
        RECT 95.745 162.025 95.915 162.195 ;
        RECT 96.205 162.025 96.375 162.195 ;
        RECT 96.665 162.025 96.835 162.195 ;
        RECT 97.125 162.025 97.295 162.195 ;
        RECT 97.585 162.025 97.755 162.195 ;
        RECT 98.045 162.025 98.215 162.195 ;
        RECT 98.505 162.025 98.675 162.195 ;
        RECT 98.965 162.025 99.135 162.195 ;
        RECT 99.425 162.025 99.595 162.195 ;
        RECT 99.885 162.025 100.055 162.195 ;
        RECT 100.345 162.025 100.515 162.195 ;
        RECT 100.805 162.025 100.975 162.195 ;
        RECT 101.265 162.025 101.435 162.195 ;
        RECT 101.725 162.025 101.895 162.195 ;
        RECT 102.185 162.025 102.355 162.195 ;
        RECT 102.645 162.025 102.815 162.195 ;
        RECT 103.105 162.025 103.275 162.195 ;
        RECT 103.565 162.025 103.735 162.195 ;
        RECT 104.025 162.025 104.195 162.195 ;
        RECT 104.485 162.025 104.655 162.195 ;
        RECT 104.945 162.025 105.115 162.195 ;
        RECT 105.405 162.025 105.575 162.195 ;
        RECT 105.865 162.025 106.035 162.195 ;
        RECT 106.325 162.025 106.495 162.195 ;
        RECT 106.785 162.025 106.955 162.195 ;
        RECT 107.245 162.025 107.415 162.195 ;
        RECT 107.705 162.025 107.875 162.195 ;
        RECT 108.165 162.025 108.335 162.195 ;
        RECT 108.625 162.025 108.795 162.195 ;
        RECT 109.085 162.025 109.255 162.195 ;
        RECT 109.545 162.025 109.715 162.195 ;
        RECT 110.005 162.025 110.175 162.195 ;
        RECT 110.465 162.025 110.635 162.195 ;
        RECT 110.925 162.025 111.095 162.195 ;
        RECT 111.385 162.025 111.555 162.195 ;
        RECT 111.845 162.025 112.015 162.195 ;
        RECT 112.305 162.025 112.475 162.195 ;
        RECT 112.765 162.025 112.935 162.195 ;
        RECT 113.225 162.025 113.395 162.195 ;
        RECT 113.685 162.025 113.855 162.195 ;
        RECT 114.145 162.025 114.315 162.195 ;
        RECT 114.605 162.025 114.775 162.195 ;
        RECT 115.065 162.025 115.235 162.195 ;
        RECT 115.525 162.025 115.695 162.195 ;
        RECT 41.925 156.585 42.095 156.755 ;
        RECT 42.385 156.585 42.555 156.755 ;
        RECT 42.845 156.585 43.015 156.755 ;
        RECT 43.305 156.585 43.475 156.755 ;
        RECT 43.765 156.585 43.935 156.755 ;
        RECT 44.225 156.585 44.395 156.755 ;
        RECT 44.685 156.585 44.855 156.755 ;
        RECT 45.145 156.585 45.315 156.755 ;
        RECT 45.605 156.585 45.775 156.755 ;
        RECT 46.065 156.585 46.235 156.755 ;
        RECT 46.525 156.585 46.695 156.755 ;
        RECT 46.985 156.585 47.155 156.755 ;
        RECT 47.445 156.585 47.615 156.755 ;
        RECT 47.905 156.585 48.075 156.755 ;
        RECT 48.365 156.585 48.535 156.755 ;
        RECT 48.825 156.585 48.995 156.755 ;
        RECT 49.285 156.585 49.455 156.755 ;
        RECT 49.745 156.585 49.915 156.755 ;
        RECT 50.205 156.585 50.375 156.755 ;
        RECT 50.665 156.585 50.835 156.755 ;
        RECT 51.125 156.585 51.295 156.755 ;
        RECT 51.585 156.585 51.755 156.755 ;
        RECT 52.045 156.585 52.215 156.755 ;
        RECT 52.505 156.585 52.675 156.755 ;
        RECT 52.965 156.585 53.135 156.755 ;
        RECT 53.425 156.585 53.595 156.755 ;
        RECT 53.885 156.585 54.055 156.755 ;
        RECT 54.345 156.585 54.515 156.755 ;
        RECT 54.805 156.585 54.975 156.755 ;
        RECT 55.265 156.585 55.435 156.755 ;
        RECT 55.725 156.585 55.895 156.755 ;
        RECT 56.185 156.585 56.355 156.755 ;
        RECT 56.645 156.585 56.815 156.755 ;
        RECT 57.105 156.585 57.275 156.755 ;
        RECT 57.565 156.585 57.735 156.755 ;
        RECT 58.025 156.585 58.195 156.755 ;
        RECT 58.485 156.585 58.655 156.755 ;
        RECT 58.945 156.585 59.115 156.755 ;
        RECT 59.405 156.585 59.575 156.755 ;
        RECT 59.865 156.585 60.035 156.755 ;
        RECT 60.325 156.585 60.495 156.755 ;
        RECT 60.785 156.585 60.955 156.755 ;
        RECT 61.245 156.585 61.415 156.755 ;
        RECT 61.705 156.585 61.875 156.755 ;
        RECT 62.165 156.585 62.335 156.755 ;
        RECT 62.625 156.585 62.795 156.755 ;
        RECT 63.085 156.585 63.255 156.755 ;
        RECT 63.545 156.585 63.715 156.755 ;
        RECT 64.005 156.585 64.175 156.755 ;
        RECT 64.465 156.585 64.635 156.755 ;
        RECT 64.925 156.585 65.095 156.755 ;
        RECT 65.385 156.585 65.555 156.755 ;
        RECT 65.845 156.585 66.015 156.755 ;
        RECT 66.305 156.585 66.475 156.755 ;
        RECT 66.765 156.585 66.935 156.755 ;
        RECT 67.225 156.585 67.395 156.755 ;
        RECT 67.685 156.585 67.855 156.755 ;
        RECT 68.145 156.585 68.315 156.755 ;
        RECT 68.605 156.585 68.775 156.755 ;
        RECT 69.065 156.585 69.235 156.755 ;
        RECT 69.525 156.585 69.695 156.755 ;
        RECT 69.985 156.585 70.155 156.755 ;
        RECT 70.445 156.585 70.615 156.755 ;
        RECT 70.905 156.585 71.075 156.755 ;
        RECT 71.365 156.585 71.535 156.755 ;
        RECT 71.825 156.585 71.995 156.755 ;
        RECT 72.285 156.585 72.455 156.755 ;
        RECT 72.745 156.585 72.915 156.755 ;
        RECT 73.205 156.585 73.375 156.755 ;
        RECT 73.665 156.585 73.835 156.755 ;
        RECT 74.125 156.585 74.295 156.755 ;
        RECT 74.585 156.585 74.755 156.755 ;
        RECT 75.045 156.585 75.215 156.755 ;
        RECT 75.505 156.585 75.675 156.755 ;
        RECT 75.965 156.585 76.135 156.755 ;
        RECT 76.425 156.585 76.595 156.755 ;
        RECT 76.885 156.585 77.055 156.755 ;
        RECT 77.345 156.585 77.515 156.755 ;
        RECT 77.805 156.585 77.975 156.755 ;
        RECT 78.265 156.585 78.435 156.755 ;
        RECT 78.725 156.585 78.895 156.755 ;
        RECT 79.185 156.585 79.355 156.755 ;
        RECT 79.645 156.585 79.815 156.755 ;
        RECT 80.105 156.585 80.275 156.755 ;
        RECT 80.565 156.585 80.735 156.755 ;
        RECT 81.025 156.585 81.195 156.755 ;
        RECT 81.485 156.585 81.655 156.755 ;
        RECT 81.945 156.585 82.115 156.755 ;
        RECT 82.405 156.585 82.575 156.755 ;
        RECT 82.865 156.585 83.035 156.755 ;
        RECT 83.325 156.585 83.495 156.755 ;
        RECT 83.785 156.585 83.955 156.755 ;
        RECT 84.245 156.585 84.415 156.755 ;
        RECT 84.705 156.585 84.875 156.755 ;
        RECT 85.165 156.585 85.335 156.755 ;
        RECT 85.625 156.585 85.795 156.755 ;
        RECT 86.085 156.585 86.255 156.755 ;
        RECT 86.545 156.585 86.715 156.755 ;
        RECT 87.005 156.585 87.175 156.755 ;
        RECT 87.465 156.585 87.635 156.755 ;
        RECT 87.925 156.585 88.095 156.755 ;
        RECT 88.385 156.585 88.555 156.755 ;
        RECT 88.845 156.585 89.015 156.755 ;
        RECT 89.305 156.585 89.475 156.755 ;
        RECT 89.765 156.585 89.935 156.755 ;
        RECT 90.225 156.585 90.395 156.755 ;
        RECT 90.685 156.585 90.855 156.755 ;
        RECT 91.145 156.585 91.315 156.755 ;
        RECT 91.605 156.585 91.775 156.755 ;
        RECT 92.065 156.585 92.235 156.755 ;
        RECT 92.525 156.585 92.695 156.755 ;
        RECT 92.985 156.585 93.155 156.755 ;
        RECT 93.445 156.585 93.615 156.755 ;
        RECT 93.905 156.585 94.075 156.755 ;
        RECT 94.365 156.585 94.535 156.755 ;
        RECT 94.825 156.585 94.995 156.755 ;
        RECT 95.285 156.585 95.455 156.755 ;
        RECT 95.745 156.585 95.915 156.755 ;
        RECT 96.205 156.585 96.375 156.755 ;
        RECT 96.665 156.585 96.835 156.755 ;
        RECT 97.125 156.585 97.295 156.755 ;
        RECT 97.585 156.585 97.755 156.755 ;
        RECT 98.045 156.585 98.215 156.755 ;
        RECT 98.505 156.585 98.675 156.755 ;
        RECT 98.965 156.585 99.135 156.755 ;
        RECT 99.425 156.585 99.595 156.755 ;
        RECT 99.885 156.585 100.055 156.755 ;
        RECT 100.345 156.585 100.515 156.755 ;
        RECT 100.805 156.585 100.975 156.755 ;
        RECT 101.265 156.585 101.435 156.755 ;
        RECT 101.725 156.585 101.895 156.755 ;
        RECT 102.185 156.585 102.355 156.755 ;
        RECT 102.645 156.585 102.815 156.755 ;
        RECT 103.105 156.585 103.275 156.755 ;
        RECT 103.565 156.585 103.735 156.755 ;
        RECT 104.025 156.585 104.195 156.755 ;
        RECT 104.485 156.585 104.655 156.755 ;
        RECT 104.945 156.585 105.115 156.755 ;
        RECT 105.405 156.585 105.575 156.755 ;
        RECT 105.865 156.585 106.035 156.755 ;
        RECT 106.325 156.585 106.495 156.755 ;
        RECT 106.785 156.585 106.955 156.755 ;
        RECT 107.245 156.585 107.415 156.755 ;
        RECT 107.705 156.585 107.875 156.755 ;
        RECT 108.165 156.585 108.335 156.755 ;
        RECT 108.625 156.585 108.795 156.755 ;
        RECT 109.085 156.585 109.255 156.755 ;
        RECT 109.545 156.585 109.715 156.755 ;
        RECT 110.005 156.585 110.175 156.755 ;
        RECT 110.465 156.585 110.635 156.755 ;
        RECT 110.925 156.585 111.095 156.755 ;
        RECT 111.385 156.585 111.555 156.755 ;
        RECT 111.845 156.585 112.015 156.755 ;
        RECT 112.305 156.585 112.475 156.755 ;
        RECT 112.765 156.585 112.935 156.755 ;
        RECT 113.225 156.585 113.395 156.755 ;
        RECT 113.685 156.585 113.855 156.755 ;
        RECT 114.145 156.585 114.315 156.755 ;
        RECT 114.605 156.585 114.775 156.755 ;
        RECT 115.065 156.585 115.235 156.755 ;
        RECT 115.525 156.585 115.695 156.755 ;
        RECT 63.940 125.590 64.110 127.470 ;
        RECT 64.530 125.590 64.700 127.470 ;
        RECT 70.170 125.590 70.340 127.470 ;
        RECT 72.050 125.590 72.220 127.470 ;
        RECT 73.930 125.590 74.100 127.470 ;
        RECT 76.650 126.770 76.860 126.980 ;
        RECT 76.650 125.480 76.860 125.690 ;
        RECT 86.600 125.590 86.770 127.470 ;
        RECT 87.190 125.590 87.360 127.470 ;
        RECT 92.830 125.590 93.000 127.470 ;
        RECT 94.710 125.590 94.880 127.470 ;
        RECT 96.590 125.590 96.760 127.470 ;
        RECT 99.310 126.770 99.520 126.980 ;
        RECT 99.310 125.480 99.520 125.690 ;
        RECT 109.260 125.590 109.430 127.470 ;
        RECT 109.850 125.590 110.020 127.470 ;
        RECT 115.490 125.590 115.660 127.470 ;
        RECT 117.370 125.590 117.540 127.470 ;
        RECT 119.250 125.590 119.420 127.470 ;
        RECT 121.970 126.770 122.180 126.980 ;
        RECT 121.970 125.480 122.180 125.690 ;
        RECT 124.280 124.705 124.470 126.690 ;
        RECT 58.155 122.545 58.325 122.715 ;
        RECT 63.940 122.500 64.110 124.380 ;
        RECT 64.530 122.500 64.700 124.380 ;
        RECT 70.170 122.500 70.340 124.380 ;
        RECT 72.050 122.500 72.220 124.380 ;
        RECT 73.930 122.500 74.100 124.380 ;
        RECT 76.650 124.195 76.860 124.405 ;
        RECT 76.650 122.910 76.860 123.120 ;
        RECT 80.815 122.545 80.985 122.715 ;
        RECT 86.600 122.500 86.770 124.380 ;
        RECT 87.190 122.500 87.360 124.380 ;
        RECT 92.830 122.500 93.000 124.380 ;
        RECT 94.710 122.500 94.880 124.380 ;
        RECT 96.590 122.500 96.760 124.380 ;
        RECT 99.310 124.195 99.520 124.405 ;
        RECT 99.310 122.910 99.520 123.120 ;
        RECT 103.475 122.545 103.645 122.715 ;
        RECT 109.260 122.500 109.430 124.380 ;
        RECT 109.850 122.500 110.020 124.380 ;
        RECT 115.490 122.500 115.660 124.380 ;
        RECT 117.370 122.500 117.540 124.380 ;
        RECT 119.250 122.500 119.420 124.380 ;
        RECT 121.970 124.195 122.180 124.405 ;
        RECT 121.970 122.910 122.180 123.120 ;
        RECT 59.470 121.700 59.640 122.080 ;
        RECT 60.870 121.700 61.040 122.080 ;
        RECT 82.130 121.700 82.300 122.080 ;
        RECT 83.530 121.700 83.700 122.080 ;
        RECT 104.790 121.700 104.960 122.080 ;
        RECT 106.190 121.700 106.360 122.080 ;
        RECT 41.280 108.250 41.450 110.130 ;
        RECT 41.870 108.250 42.040 110.130 ;
        RECT 47.510 108.250 47.680 110.130 ;
        RECT 49.390 108.250 49.560 110.130 ;
        RECT 51.270 108.250 51.440 110.130 ;
        RECT 53.990 109.430 54.200 109.640 ;
        RECT 53.990 108.140 54.200 108.350 ;
        RECT 63.940 108.250 64.110 110.130 ;
        RECT 64.530 108.250 64.700 110.130 ;
        RECT 70.170 108.250 70.340 110.130 ;
        RECT 72.050 108.250 72.220 110.130 ;
        RECT 73.930 108.250 74.100 110.130 ;
        RECT 76.650 109.430 76.860 109.640 ;
        RECT 76.650 108.140 76.860 108.350 ;
        RECT 86.600 108.250 86.770 110.130 ;
        RECT 87.190 108.250 87.360 110.130 ;
        RECT 92.830 108.250 93.000 110.130 ;
        RECT 94.710 108.250 94.880 110.130 ;
        RECT 96.590 108.250 96.760 110.130 ;
        RECT 99.310 109.430 99.520 109.640 ;
        RECT 99.310 108.140 99.520 108.350 ;
        RECT 109.260 108.250 109.430 110.130 ;
        RECT 109.850 108.250 110.020 110.130 ;
        RECT 115.490 108.250 115.660 110.130 ;
        RECT 117.370 108.250 117.540 110.130 ;
        RECT 119.250 108.250 119.420 110.130 ;
        RECT 121.970 109.430 122.180 109.640 ;
        RECT 121.970 108.140 122.180 108.350 ;
        RECT 35.495 105.205 35.665 105.375 ;
        RECT 41.280 105.160 41.450 107.040 ;
        RECT 41.870 105.160 42.040 107.040 ;
        RECT 47.510 105.160 47.680 107.040 ;
        RECT 49.390 105.160 49.560 107.040 ;
        RECT 51.270 105.160 51.440 107.040 ;
        RECT 53.990 106.855 54.200 107.065 ;
        RECT 53.990 105.570 54.200 105.780 ;
        RECT 58.155 105.205 58.325 105.375 ;
        RECT 63.940 105.160 64.110 107.040 ;
        RECT 64.530 105.160 64.700 107.040 ;
        RECT 70.170 105.160 70.340 107.040 ;
        RECT 72.050 105.160 72.220 107.040 ;
        RECT 73.930 105.160 74.100 107.040 ;
        RECT 76.650 106.855 76.860 107.065 ;
        RECT 76.650 105.570 76.860 105.780 ;
        RECT 80.815 105.205 80.985 105.375 ;
        RECT 86.600 105.160 86.770 107.040 ;
        RECT 87.190 105.160 87.360 107.040 ;
        RECT 92.830 105.160 93.000 107.040 ;
        RECT 94.710 105.160 94.880 107.040 ;
        RECT 96.590 105.160 96.760 107.040 ;
        RECT 99.310 106.855 99.520 107.065 ;
        RECT 99.310 105.570 99.520 105.780 ;
        RECT 103.475 105.205 103.645 105.375 ;
        RECT 109.260 105.160 109.430 107.040 ;
        RECT 109.850 105.160 110.020 107.040 ;
        RECT 115.490 105.160 115.660 107.040 ;
        RECT 117.370 105.160 117.540 107.040 ;
        RECT 119.250 105.160 119.420 107.040 ;
        RECT 121.970 106.855 122.180 107.065 ;
        RECT 121.970 105.570 122.180 105.780 ;
        RECT 36.810 104.360 36.980 104.740 ;
        RECT 38.210 104.360 38.380 104.740 ;
        RECT 59.470 104.360 59.640 104.740 ;
        RECT 60.870 104.360 61.040 104.740 ;
        RECT 82.130 104.360 82.300 104.740 ;
        RECT 83.530 104.360 83.700 104.740 ;
        RECT 104.790 104.360 104.960 104.740 ;
        RECT 106.190 104.360 106.360 104.740 ;
        RECT 41.280 90.910 41.450 92.790 ;
        RECT 41.870 90.910 42.040 92.790 ;
        RECT 47.510 90.910 47.680 92.790 ;
        RECT 49.390 90.910 49.560 92.790 ;
        RECT 51.270 90.910 51.440 92.790 ;
        RECT 53.990 92.090 54.200 92.300 ;
        RECT 53.990 90.800 54.200 91.010 ;
        RECT 63.940 90.910 64.110 92.790 ;
        RECT 64.530 90.910 64.700 92.790 ;
        RECT 70.170 90.910 70.340 92.790 ;
        RECT 72.050 90.910 72.220 92.790 ;
        RECT 73.930 90.910 74.100 92.790 ;
        RECT 76.650 92.090 76.860 92.300 ;
        RECT 76.650 90.800 76.860 91.010 ;
        RECT 86.600 90.910 86.770 92.790 ;
        RECT 87.190 90.910 87.360 92.790 ;
        RECT 92.830 90.910 93.000 92.790 ;
        RECT 94.710 90.910 94.880 92.790 ;
        RECT 96.590 90.910 96.760 92.790 ;
        RECT 99.310 92.090 99.520 92.300 ;
        RECT 99.310 90.800 99.520 91.010 ;
        RECT 109.260 90.910 109.430 92.790 ;
        RECT 109.850 90.910 110.020 92.790 ;
        RECT 115.490 90.910 115.660 92.790 ;
        RECT 117.370 90.910 117.540 92.790 ;
        RECT 119.250 90.910 119.420 92.790 ;
        RECT 121.970 92.090 122.180 92.300 ;
        RECT 121.970 90.800 122.180 91.010 ;
        RECT 35.495 87.865 35.665 88.035 ;
        RECT 41.280 87.820 41.450 89.700 ;
        RECT 41.870 87.820 42.040 89.700 ;
        RECT 47.510 87.820 47.680 89.700 ;
        RECT 49.390 87.820 49.560 89.700 ;
        RECT 51.270 87.820 51.440 89.700 ;
        RECT 53.990 89.515 54.200 89.725 ;
        RECT 53.990 88.230 54.200 88.440 ;
        RECT 58.155 87.865 58.325 88.035 ;
        RECT 63.940 87.820 64.110 89.700 ;
        RECT 64.530 87.820 64.700 89.700 ;
        RECT 70.170 87.820 70.340 89.700 ;
        RECT 72.050 87.820 72.220 89.700 ;
        RECT 73.930 87.820 74.100 89.700 ;
        RECT 76.650 89.515 76.860 89.725 ;
        RECT 76.650 88.230 76.860 88.440 ;
        RECT 80.815 87.865 80.985 88.035 ;
        RECT 86.600 87.820 86.770 89.700 ;
        RECT 87.190 87.820 87.360 89.700 ;
        RECT 92.830 87.820 93.000 89.700 ;
        RECT 94.710 87.820 94.880 89.700 ;
        RECT 96.590 87.820 96.760 89.700 ;
        RECT 99.310 89.515 99.520 89.725 ;
        RECT 99.310 88.230 99.520 88.440 ;
        RECT 103.475 87.865 103.645 88.035 ;
        RECT 109.260 87.820 109.430 89.700 ;
        RECT 109.850 87.820 110.020 89.700 ;
        RECT 115.490 87.820 115.660 89.700 ;
        RECT 117.370 87.820 117.540 89.700 ;
        RECT 119.250 87.820 119.420 89.700 ;
        RECT 121.970 89.515 122.180 89.725 ;
        RECT 121.970 88.230 122.180 88.440 ;
        RECT 36.810 87.020 36.980 87.400 ;
        RECT 38.210 87.020 38.380 87.400 ;
        RECT 59.470 87.020 59.640 87.400 ;
        RECT 60.870 87.020 61.040 87.400 ;
        RECT 82.130 87.020 82.300 87.400 ;
        RECT 83.530 87.020 83.700 87.400 ;
        RECT 104.790 87.020 104.960 87.400 ;
        RECT 106.190 87.020 106.360 87.400 ;
        RECT 41.280 73.570 41.450 75.450 ;
        RECT 41.870 73.570 42.040 75.450 ;
        RECT 47.510 73.570 47.680 75.450 ;
        RECT 49.390 73.570 49.560 75.450 ;
        RECT 51.270 73.570 51.440 75.450 ;
        RECT 53.990 74.750 54.200 74.960 ;
        RECT 53.990 73.460 54.200 73.670 ;
        RECT 63.940 73.570 64.110 75.450 ;
        RECT 64.530 73.570 64.700 75.450 ;
        RECT 70.170 73.570 70.340 75.450 ;
        RECT 72.050 73.570 72.220 75.450 ;
        RECT 73.930 73.570 74.100 75.450 ;
        RECT 76.650 74.750 76.860 74.960 ;
        RECT 76.650 73.460 76.860 73.670 ;
        RECT 86.600 73.570 86.770 75.450 ;
        RECT 87.190 73.570 87.360 75.450 ;
        RECT 92.830 73.570 93.000 75.450 ;
        RECT 94.710 73.570 94.880 75.450 ;
        RECT 96.590 73.570 96.760 75.450 ;
        RECT 99.310 74.750 99.520 74.960 ;
        RECT 99.310 73.460 99.520 73.670 ;
        RECT 109.260 73.570 109.430 75.450 ;
        RECT 109.850 73.570 110.020 75.450 ;
        RECT 115.490 73.570 115.660 75.450 ;
        RECT 117.370 73.570 117.540 75.450 ;
        RECT 119.250 73.570 119.420 75.450 ;
        RECT 121.970 74.750 122.180 74.960 ;
        RECT 121.970 73.460 122.180 73.670 ;
        RECT 35.495 70.525 35.665 70.695 ;
        RECT 41.280 70.480 41.450 72.360 ;
        RECT 41.870 70.480 42.040 72.360 ;
        RECT 47.510 70.480 47.680 72.360 ;
        RECT 49.390 70.480 49.560 72.360 ;
        RECT 51.270 70.480 51.440 72.360 ;
        RECT 53.990 72.175 54.200 72.385 ;
        RECT 53.990 70.890 54.200 71.100 ;
        RECT 58.155 70.525 58.325 70.695 ;
        RECT 63.940 70.480 64.110 72.360 ;
        RECT 64.530 70.480 64.700 72.360 ;
        RECT 70.170 70.480 70.340 72.360 ;
        RECT 72.050 70.480 72.220 72.360 ;
        RECT 73.930 70.480 74.100 72.360 ;
        RECT 76.650 72.175 76.860 72.385 ;
        RECT 76.650 70.890 76.860 71.100 ;
        RECT 80.815 70.525 80.985 70.695 ;
        RECT 86.600 70.480 86.770 72.360 ;
        RECT 87.190 70.480 87.360 72.360 ;
        RECT 92.830 70.480 93.000 72.360 ;
        RECT 94.710 70.480 94.880 72.360 ;
        RECT 96.590 70.480 96.760 72.360 ;
        RECT 99.310 72.175 99.520 72.385 ;
        RECT 99.310 70.890 99.520 71.100 ;
        RECT 103.475 70.525 103.645 70.695 ;
        RECT 109.260 70.480 109.430 72.360 ;
        RECT 109.850 70.480 110.020 72.360 ;
        RECT 115.490 70.480 115.660 72.360 ;
        RECT 117.370 70.480 117.540 72.360 ;
        RECT 119.250 70.480 119.420 72.360 ;
        RECT 121.970 72.175 122.180 72.385 ;
        RECT 121.970 70.890 122.180 71.100 ;
        RECT 36.810 69.680 36.980 70.060 ;
        RECT 38.210 69.680 38.380 70.060 ;
        RECT 59.470 69.680 59.640 70.060 ;
        RECT 60.870 69.680 61.040 70.060 ;
        RECT 82.130 69.680 82.300 70.060 ;
        RECT 83.530 69.680 83.700 70.060 ;
        RECT 104.790 69.680 104.960 70.060 ;
        RECT 106.190 69.680 106.360 70.060 ;
        RECT 41.280 55.570 41.450 57.450 ;
        RECT 41.870 55.570 42.040 57.450 ;
        RECT 47.510 55.570 47.680 57.450 ;
        RECT 49.390 55.570 49.560 57.450 ;
        RECT 51.270 55.570 51.440 57.450 ;
        RECT 53.990 56.750 54.200 56.960 ;
        RECT 53.990 55.460 54.200 55.670 ;
        RECT 63.940 55.570 64.110 57.450 ;
        RECT 64.530 55.570 64.700 57.450 ;
        RECT 70.170 55.570 70.340 57.450 ;
        RECT 72.050 55.570 72.220 57.450 ;
        RECT 73.930 55.570 74.100 57.450 ;
        RECT 76.650 56.750 76.860 56.960 ;
        RECT 76.650 55.460 76.860 55.670 ;
        RECT 86.600 55.570 86.770 57.450 ;
        RECT 87.190 55.570 87.360 57.450 ;
        RECT 92.830 55.570 93.000 57.450 ;
        RECT 94.710 55.570 94.880 57.450 ;
        RECT 96.590 55.570 96.760 57.450 ;
        RECT 99.310 56.750 99.520 56.960 ;
        RECT 99.310 55.460 99.520 55.670 ;
        RECT 109.260 55.570 109.430 57.450 ;
        RECT 109.850 55.570 110.020 57.450 ;
        RECT 115.490 55.570 115.660 57.450 ;
        RECT 117.370 55.570 117.540 57.450 ;
        RECT 119.250 55.570 119.420 57.450 ;
        RECT 121.970 56.750 122.180 56.960 ;
        RECT 121.970 55.460 122.180 55.670 ;
        RECT 41.280 52.480 41.450 54.360 ;
        RECT 41.870 52.480 42.040 54.360 ;
        RECT 47.510 52.480 47.680 54.360 ;
        RECT 49.390 52.480 49.560 54.360 ;
        RECT 51.270 52.480 51.440 54.360 ;
        RECT 53.990 54.175 54.200 54.385 ;
        RECT 53.990 52.890 54.200 53.100 ;
        RECT 63.940 52.480 64.110 54.360 ;
        RECT 64.530 52.480 64.700 54.360 ;
        RECT 70.170 52.480 70.340 54.360 ;
        RECT 72.050 52.480 72.220 54.360 ;
        RECT 73.930 52.480 74.100 54.360 ;
        RECT 76.650 54.175 76.860 54.385 ;
        RECT 76.650 52.890 76.860 53.100 ;
        RECT 86.600 52.480 86.770 54.360 ;
        RECT 87.190 52.480 87.360 54.360 ;
        RECT 92.830 52.480 93.000 54.360 ;
        RECT 94.710 52.480 94.880 54.360 ;
        RECT 96.590 52.480 96.760 54.360 ;
        RECT 99.310 54.175 99.520 54.385 ;
        RECT 99.310 52.890 99.520 53.100 ;
        RECT 109.260 52.480 109.430 54.360 ;
        RECT 109.850 52.480 110.020 54.360 ;
        RECT 115.490 52.480 115.660 54.360 ;
        RECT 117.370 52.480 117.540 54.360 ;
        RECT 119.250 52.480 119.420 54.360 ;
        RECT 121.970 54.175 122.180 54.385 ;
        RECT 121.970 52.890 122.180 53.100 ;
      LAYER met1 ;
        RECT 41.780 183.630 116.620 184.110 ;
        RECT 41.780 178.190 116.620 178.670 ;
        RECT 41.780 172.750 116.620 173.230 ;
        RECT 41.780 167.310 116.620 167.790 ;
        RECT 41.780 161.870 116.620 162.350 ;
        RECT 41.780 156.430 116.620 156.910 ;
        RECT 63.910 127.500 64.140 127.530 ;
        RECT 64.500 127.500 64.730 127.530 ;
        RECT 63.910 126.900 64.730 127.500 ;
        RECT 70.060 126.930 70.660 127.530 ;
        RECT 71.940 126.930 72.540 127.530 ;
        RECT 73.820 126.930 74.420 127.530 ;
        RECT 86.570 127.500 86.800 127.530 ;
        RECT 87.160 127.500 87.390 127.530 ;
        RECT 75.630 127.020 75.890 127.340 ;
        RECT 76.660 127.070 76.850 127.100 ;
        RECT 75.665 126.970 75.890 127.020 ;
        RECT 76.620 126.970 76.890 127.070 ;
        RECT 63.910 125.780 64.140 126.900 ;
        RECT 64.500 125.780 64.730 126.900 ;
        RECT 63.910 125.530 64.730 125.780 ;
        RECT 70.140 125.775 70.370 126.930 ;
        RECT 72.020 125.785 72.250 126.930 ;
        RECT 73.900 125.785 74.130 126.930 ;
        RECT 70.055 125.530 70.370 125.775 ;
        RECT 71.925 125.530 72.250 125.785 ;
        RECT 73.805 125.530 74.130 125.785 ;
        RECT 75.665 126.780 76.890 126.970 ;
        RECT 75.665 125.680 75.855 126.780 ;
        RECT 76.620 126.690 76.890 126.780 ;
        RECT 86.570 126.900 87.390 127.500 ;
        RECT 92.720 126.930 93.320 127.530 ;
        RECT 94.600 126.930 95.200 127.530 ;
        RECT 96.480 126.930 97.080 127.530 ;
        RECT 109.230 127.500 109.460 127.530 ;
        RECT 109.820 127.500 110.050 127.530 ;
        RECT 98.290 127.020 98.550 127.340 ;
        RECT 99.320 127.070 99.510 127.100 ;
        RECT 98.325 126.970 98.550 127.020 ;
        RECT 99.280 126.970 99.550 127.070 ;
        RECT 76.660 125.780 76.850 125.810 ;
        RECT 86.570 125.780 86.800 126.900 ;
        RECT 87.160 125.780 87.390 126.900 ;
        RECT 76.620 125.680 76.890 125.780 ;
        RECT 64.030 124.440 64.595 125.530 ;
        RECT 70.055 124.440 70.245 125.530 ;
        RECT 71.925 124.440 72.115 125.530 ;
        RECT 73.805 124.440 73.995 125.530 ;
        RECT 75.665 125.490 76.890 125.680 ;
        RECT 86.570 125.530 87.390 125.780 ;
        RECT 92.800 125.775 93.030 126.930 ;
        RECT 94.680 125.785 94.910 126.930 ;
        RECT 96.560 125.785 96.790 126.930 ;
        RECT 92.715 125.530 93.030 125.775 ;
        RECT 94.585 125.530 94.910 125.785 ;
        RECT 96.465 125.530 96.790 125.785 ;
        RECT 98.325 126.780 99.550 126.970 ;
        RECT 98.325 125.680 98.515 126.780 ;
        RECT 99.280 126.690 99.550 126.780 ;
        RECT 109.230 126.900 110.050 127.500 ;
        RECT 115.380 126.930 115.980 127.530 ;
        RECT 117.260 126.930 117.860 127.530 ;
        RECT 119.140 126.930 119.740 127.530 ;
        RECT 120.950 127.020 121.210 127.340 ;
        RECT 121.980 127.070 122.170 127.100 ;
        RECT 120.985 126.970 121.210 127.020 ;
        RECT 121.940 126.970 122.210 127.070 ;
        RECT 99.320 125.780 99.510 125.810 ;
        RECT 109.230 125.780 109.460 126.900 ;
        RECT 109.820 125.780 110.050 126.900 ;
        RECT 99.280 125.680 99.550 125.780 ;
        RECT 63.910 124.200 64.730 124.440 ;
        RECT 70.055 124.200 70.370 124.440 ;
        RECT 71.925 124.200 72.250 124.440 ;
        RECT 58.450 122.745 61.435 122.875 ;
        RECT 58.095 122.685 61.435 122.745 ;
        RECT 58.095 122.535 58.650 122.685 ;
        RECT 58.095 122.515 58.385 122.535 ;
        RECT 59.645 122.140 59.835 122.685 ;
        RECT 61.245 122.580 61.435 122.685 ;
        RECT 63.910 122.680 64.140 124.200 ;
        RECT 64.500 122.680 64.730 124.200 ;
        RECT 61.245 122.425 62.250 122.580 ;
        RECT 63.910 122.490 64.730 122.680 ;
        RECT 63.910 122.440 64.140 122.490 ;
        RECT 64.500 122.440 64.730 122.490 ;
        RECT 70.140 122.440 70.370 124.200 ;
        RECT 72.020 122.440 72.250 124.200 ;
        RECT 73.805 124.195 74.130 124.440 ;
        RECT 73.900 122.440 74.130 124.195 ;
        RECT 75.665 124.395 75.855 125.490 ;
        RECT 76.620 125.400 76.890 125.490 ;
        RECT 76.660 124.495 76.850 124.525 ;
        RECT 76.620 124.395 76.890 124.495 ;
        RECT 86.690 124.440 87.255 125.530 ;
        RECT 92.715 124.440 92.905 125.530 ;
        RECT 94.585 124.440 94.775 125.530 ;
        RECT 96.465 124.440 96.655 125.530 ;
        RECT 98.325 125.490 99.550 125.680 ;
        RECT 109.230 125.530 110.050 125.780 ;
        RECT 115.460 125.775 115.690 126.930 ;
        RECT 117.340 125.785 117.570 126.930 ;
        RECT 119.220 125.785 119.450 126.930 ;
        RECT 115.375 125.530 115.690 125.775 ;
        RECT 117.245 125.530 117.570 125.785 ;
        RECT 119.125 125.530 119.450 125.785 ;
        RECT 120.985 126.780 122.210 126.970 ;
        RECT 120.985 125.680 121.175 126.780 ;
        RECT 121.940 126.690 122.210 126.780 ;
        RECT 121.980 125.780 122.170 125.810 ;
        RECT 121.940 125.680 122.210 125.780 ;
        RECT 75.665 124.205 76.890 124.395 ;
        RECT 75.665 123.110 75.855 124.205 ;
        RECT 76.620 124.115 76.890 124.205 ;
        RECT 86.570 124.200 87.390 124.440 ;
        RECT 92.715 124.200 93.030 124.440 ;
        RECT 94.585 124.200 94.910 124.440 ;
        RECT 76.660 123.210 76.850 123.245 ;
        RECT 76.620 123.110 76.890 123.210 ;
        RECT 75.665 122.920 76.890 123.110 ;
        RECT 76.620 122.830 76.890 122.920 ;
        RECT 81.110 122.745 84.095 122.875 ;
        RECT 80.755 122.685 84.095 122.745 ;
        RECT 80.755 122.535 81.310 122.685 ;
        RECT 80.755 122.515 81.045 122.535 ;
        RECT 59.440 121.950 59.835 122.140 ;
        RECT 60.840 122.090 61.070 122.140 ;
        RECT 61.250 122.090 62.250 122.425 ;
        RECT 82.305 122.140 82.495 122.685 ;
        RECT 83.905 122.580 84.095 122.685 ;
        RECT 86.570 122.680 86.800 124.200 ;
        RECT 87.160 122.680 87.390 124.200 ;
        RECT 83.905 122.425 84.910 122.580 ;
        RECT 86.570 122.490 87.390 122.680 ;
        RECT 86.570 122.440 86.800 122.490 ;
        RECT 87.160 122.440 87.390 122.490 ;
        RECT 92.800 122.440 93.030 124.200 ;
        RECT 94.680 122.440 94.910 124.200 ;
        RECT 96.465 124.195 96.790 124.440 ;
        RECT 96.560 122.440 96.790 124.195 ;
        RECT 98.325 124.395 98.515 125.490 ;
        RECT 99.280 125.400 99.550 125.490 ;
        RECT 99.320 124.495 99.510 124.525 ;
        RECT 99.280 124.395 99.550 124.495 ;
        RECT 109.350 124.440 109.915 125.530 ;
        RECT 115.375 124.440 115.565 125.530 ;
        RECT 117.245 124.440 117.435 125.530 ;
        RECT 119.125 124.440 119.315 125.530 ;
        RECT 120.985 125.490 122.210 125.680 ;
        RECT 98.325 124.205 99.550 124.395 ;
        RECT 98.325 123.110 98.515 124.205 ;
        RECT 99.280 124.115 99.550 124.205 ;
        RECT 109.230 124.200 110.050 124.440 ;
        RECT 115.375 124.200 115.690 124.440 ;
        RECT 117.245 124.200 117.570 124.440 ;
        RECT 99.320 123.210 99.510 123.245 ;
        RECT 99.280 123.110 99.550 123.210 ;
        RECT 98.325 122.920 99.550 123.110 ;
        RECT 99.280 122.830 99.550 122.920 ;
        RECT 103.770 122.745 106.755 122.875 ;
        RECT 103.415 122.685 106.755 122.745 ;
        RECT 103.415 122.535 103.970 122.685 ;
        RECT 103.415 122.515 103.705 122.535 ;
        RECT 59.440 121.640 59.670 121.950 ;
        RECT 60.840 121.900 62.250 122.090 ;
        RECT 60.840 121.640 61.070 121.900 ;
        RECT 61.250 121.580 62.250 121.900 ;
        RECT 82.100 121.950 82.495 122.140 ;
        RECT 83.500 122.090 83.730 122.140 ;
        RECT 83.910 122.090 84.910 122.425 ;
        RECT 104.965 122.140 105.155 122.685 ;
        RECT 106.565 122.580 106.755 122.685 ;
        RECT 109.230 122.680 109.460 124.200 ;
        RECT 109.820 122.680 110.050 124.200 ;
        RECT 106.565 122.425 107.570 122.580 ;
        RECT 109.230 122.490 110.050 122.680 ;
        RECT 109.230 122.440 109.460 122.490 ;
        RECT 109.820 122.440 110.050 122.490 ;
        RECT 115.460 122.440 115.690 124.200 ;
        RECT 117.340 122.440 117.570 124.200 ;
        RECT 119.125 124.195 119.450 124.440 ;
        RECT 119.220 122.440 119.450 124.195 ;
        RECT 120.985 124.395 121.175 125.490 ;
        RECT 121.940 125.400 122.210 125.490 ;
        RECT 124.200 124.590 124.550 126.810 ;
        RECT 121.980 124.495 122.170 124.525 ;
        RECT 121.940 124.395 122.210 124.495 ;
        RECT 120.985 124.205 122.210 124.395 ;
        RECT 120.985 123.110 121.175 124.205 ;
        RECT 121.940 124.115 122.210 124.205 ;
        RECT 121.980 123.210 122.170 123.245 ;
        RECT 121.940 123.110 122.210 123.210 ;
        RECT 120.985 122.920 122.210 123.110 ;
        RECT 121.940 122.830 122.210 122.920 ;
        RECT 82.100 121.640 82.330 121.950 ;
        RECT 83.500 121.900 84.910 122.090 ;
        RECT 83.500 121.640 83.730 121.900 ;
        RECT 83.910 121.580 84.910 121.900 ;
        RECT 104.760 121.950 105.155 122.140 ;
        RECT 106.160 122.090 106.390 122.140 ;
        RECT 106.570 122.090 107.570 122.425 ;
        RECT 104.760 121.640 104.990 121.950 ;
        RECT 106.160 121.900 107.570 122.090 ;
        RECT 106.160 121.640 106.390 121.900 ;
        RECT 106.570 121.580 107.570 121.900 ;
        RECT 41.250 110.160 41.480 110.190 ;
        RECT 41.840 110.160 42.070 110.190 ;
        RECT 41.250 109.560 42.070 110.160 ;
        RECT 47.400 109.590 48.000 110.190 ;
        RECT 49.280 109.590 49.880 110.190 ;
        RECT 51.160 109.590 51.760 110.190 ;
        RECT 63.910 110.160 64.140 110.190 ;
        RECT 64.500 110.160 64.730 110.190 ;
        RECT 52.970 109.680 53.230 110.000 ;
        RECT 54.000 109.730 54.190 109.760 ;
        RECT 53.005 109.630 53.230 109.680 ;
        RECT 53.960 109.630 54.230 109.730 ;
        RECT 41.250 108.440 41.480 109.560 ;
        RECT 41.840 108.440 42.070 109.560 ;
        RECT 41.250 108.190 42.070 108.440 ;
        RECT 47.480 108.435 47.710 109.590 ;
        RECT 49.360 108.445 49.590 109.590 ;
        RECT 51.240 108.445 51.470 109.590 ;
        RECT 47.395 108.190 47.710 108.435 ;
        RECT 49.265 108.190 49.590 108.445 ;
        RECT 51.145 108.190 51.470 108.445 ;
        RECT 53.005 109.440 54.230 109.630 ;
        RECT 53.005 108.340 53.195 109.440 ;
        RECT 53.960 109.350 54.230 109.440 ;
        RECT 63.910 109.560 64.730 110.160 ;
        RECT 70.060 109.590 70.660 110.190 ;
        RECT 71.940 109.590 72.540 110.190 ;
        RECT 73.820 109.590 74.420 110.190 ;
        RECT 86.570 110.160 86.800 110.190 ;
        RECT 87.160 110.160 87.390 110.190 ;
        RECT 75.630 109.680 75.890 110.000 ;
        RECT 76.660 109.730 76.850 109.760 ;
        RECT 75.665 109.630 75.890 109.680 ;
        RECT 76.620 109.630 76.890 109.730 ;
        RECT 54.000 108.440 54.190 108.470 ;
        RECT 63.910 108.440 64.140 109.560 ;
        RECT 64.500 108.440 64.730 109.560 ;
        RECT 53.960 108.340 54.230 108.440 ;
        RECT 41.370 107.100 41.935 108.190 ;
        RECT 47.395 107.100 47.585 108.190 ;
        RECT 49.265 107.100 49.455 108.190 ;
        RECT 51.145 107.100 51.335 108.190 ;
        RECT 53.005 108.150 54.230 108.340 ;
        RECT 63.910 108.190 64.730 108.440 ;
        RECT 70.140 108.435 70.370 109.590 ;
        RECT 72.020 108.445 72.250 109.590 ;
        RECT 73.900 108.445 74.130 109.590 ;
        RECT 70.055 108.190 70.370 108.435 ;
        RECT 71.925 108.190 72.250 108.445 ;
        RECT 73.805 108.190 74.130 108.445 ;
        RECT 75.665 109.440 76.890 109.630 ;
        RECT 75.665 108.340 75.855 109.440 ;
        RECT 76.620 109.350 76.890 109.440 ;
        RECT 86.570 109.560 87.390 110.160 ;
        RECT 92.720 109.590 93.320 110.190 ;
        RECT 94.600 109.590 95.200 110.190 ;
        RECT 96.480 109.590 97.080 110.190 ;
        RECT 109.230 110.160 109.460 110.190 ;
        RECT 109.820 110.160 110.050 110.190 ;
        RECT 98.290 109.680 98.550 110.000 ;
        RECT 99.320 109.730 99.510 109.760 ;
        RECT 98.325 109.630 98.550 109.680 ;
        RECT 99.280 109.630 99.550 109.730 ;
        RECT 76.660 108.440 76.850 108.470 ;
        RECT 86.570 108.440 86.800 109.560 ;
        RECT 87.160 108.440 87.390 109.560 ;
        RECT 76.620 108.340 76.890 108.440 ;
        RECT 41.250 106.860 42.070 107.100 ;
        RECT 47.395 106.860 47.710 107.100 ;
        RECT 49.265 106.860 49.590 107.100 ;
        RECT 35.790 105.405 38.775 105.535 ;
        RECT 35.435 105.345 38.775 105.405 ;
        RECT 35.435 105.195 35.990 105.345 ;
        RECT 35.435 105.175 35.725 105.195 ;
        RECT 36.985 104.800 37.175 105.345 ;
        RECT 38.585 105.240 38.775 105.345 ;
        RECT 41.250 105.340 41.480 106.860 ;
        RECT 41.840 105.340 42.070 106.860 ;
        RECT 38.585 105.085 39.590 105.240 ;
        RECT 41.250 105.150 42.070 105.340 ;
        RECT 41.250 105.100 41.480 105.150 ;
        RECT 41.840 105.100 42.070 105.150 ;
        RECT 47.480 105.100 47.710 106.860 ;
        RECT 49.360 105.100 49.590 106.860 ;
        RECT 51.145 106.855 51.470 107.100 ;
        RECT 51.240 105.100 51.470 106.855 ;
        RECT 53.005 107.055 53.195 108.150 ;
        RECT 53.960 108.060 54.230 108.150 ;
        RECT 54.000 107.155 54.190 107.185 ;
        RECT 53.960 107.055 54.230 107.155 ;
        RECT 64.030 107.100 64.595 108.190 ;
        RECT 70.055 107.100 70.245 108.190 ;
        RECT 71.925 107.100 72.115 108.190 ;
        RECT 73.805 107.100 73.995 108.190 ;
        RECT 75.665 108.150 76.890 108.340 ;
        RECT 86.570 108.190 87.390 108.440 ;
        RECT 92.800 108.435 93.030 109.590 ;
        RECT 94.680 108.445 94.910 109.590 ;
        RECT 96.560 108.445 96.790 109.590 ;
        RECT 92.715 108.190 93.030 108.435 ;
        RECT 94.585 108.190 94.910 108.445 ;
        RECT 96.465 108.190 96.790 108.445 ;
        RECT 98.325 109.440 99.550 109.630 ;
        RECT 98.325 108.340 98.515 109.440 ;
        RECT 99.280 109.350 99.550 109.440 ;
        RECT 109.230 109.560 110.050 110.160 ;
        RECT 115.380 109.590 115.980 110.190 ;
        RECT 117.260 109.590 117.860 110.190 ;
        RECT 119.140 109.590 119.740 110.190 ;
        RECT 120.950 109.680 121.210 110.000 ;
        RECT 121.980 109.730 122.170 109.760 ;
        RECT 120.985 109.630 121.210 109.680 ;
        RECT 121.940 109.630 122.210 109.730 ;
        RECT 99.320 108.440 99.510 108.470 ;
        RECT 109.230 108.440 109.460 109.560 ;
        RECT 109.820 108.440 110.050 109.560 ;
        RECT 99.280 108.340 99.550 108.440 ;
        RECT 53.005 106.865 54.230 107.055 ;
        RECT 53.005 105.770 53.195 106.865 ;
        RECT 53.960 106.775 54.230 106.865 ;
        RECT 63.910 106.860 64.730 107.100 ;
        RECT 70.055 106.860 70.370 107.100 ;
        RECT 71.925 106.860 72.250 107.100 ;
        RECT 54.000 105.870 54.190 105.905 ;
        RECT 53.960 105.770 54.230 105.870 ;
        RECT 53.005 105.580 54.230 105.770 ;
        RECT 53.960 105.490 54.230 105.580 ;
        RECT 58.450 105.405 61.435 105.535 ;
        RECT 58.095 105.345 61.435 105.405 ;
        RECT 58.095 105.195 58.650 105.345 ;
        RECT 58.095 105.175 58.385 105.195 ;
        RECT 36.780 104.610 37.175 104.800 ;
        RECT 38.180 104.750 38.410 104.800 ;
        RECT 38.590 104.750 39.590 105.085 ;
        RECT 59.645 104.800 59.835 105.345 ;
        RECT 61.245 105.240 61.435 105.345 ;
        RECT 63.910 105.340 64.140 106.860 ;
        RECT 64.500 105.340 64.730 106.860 ;
        RECT 61.245 105.085 62.250 105.240 ;
        RECT 63.910 105.150 64.730 105.340 ;
        RECT 63.910 105.100 64.140 105.150 ;
        RECT 64.500 105.100 64.730 105.150 ;
        RECT 70.140 105.100 70.370 106.860 ;
        RECT 72.020 105.100 72.250 106.860 ;
        RECT 73.805 106.855 74.130 107.100 ;
        RECT 73.900 105.100 74.130 106.855 ;
        RECT 75.665 107.055 75.855 108.150 ;
        RECT 76.620 108.060 76.890 108.150 ;
        RECT 76.660 107.155 76.850 107.185 ;
        RECT 76.620 107.055 76.890 107.155 ;
        RECT 86.690 107.100 87.255 108.190 ;
        RECT 92.715 107.100 92.905 108.190 ;
        RECT 94.585 107.100 94.775 108.190 ;
        RECT 96.465 107.100 96.655 108.190 ;
        RECT 98.325 108.150 99.550 108.340 ;
        RECT 109.230 108.190 110.050 108.440 ;
        RECT 115.460 108.435 115.690 109.590 ;
        RECT 117.340 108.445 117.570 109.590 ;
        RECT 119.220 108.445 119.450 109.590 ;
        RECT 115.375 108.190 115.690 108.435 ;
        RECT 117.245 108.190 117.570 108.445 ;
        RECT 119.125 108.190 119.450 108.445 ;
        RECT 120.985 109.440 122.210 109.630 ;
        RECT 120.985 108.340 121.175 109.440 ;
        RECT 121.940 109.350 122.210 109.440 ;
        RECT 121.980 108.440 122.170 108.470 ;
        RECT 121.940 108.340 122.210 108.440 ;
        RECT 75.665 106.865 76.890 107.055 ;
        RECT 75.665 105.770 75.855 106.865 ;
        RECT 76.620 106.775 76.890 106.865 ;
        RECT 86.570 106.860 87.390 107.100 ;
        RECT 92.715 106.860 93.030 107.100 ;
        RECT 94.585 106.860 94.910 107.100 ;
        RECT 76.660 105.870 76.850 105.905 ;
        RECT 76.620 105.770 76.890 105.870 ;
        RECT 75.665 105.580 76.890 105.770 ;
        RECT 76.620 105.490 76.890 105.580 ;
        RECT 81.110 105.405 84.095 105.535 ;
        RECT 80.755 105.345 84.095 105.405 ;
        RECT 80.755 105.195 81.310 105.345 ;
        RECT 80.755 105.175 81.045 105.195 ;
        RECT 36.780 104.300 37.010 104.610 ;
        RECT 38.180 104.560 39.590 104.750 ;
        RECT 38.180 104.300 38.410 104.560 ;
        RECT 38.590 104.240 39.590 104.560 ;
        RECT 59.440 104.610 59.835 104.800 ;
        RECT 60.840 104.750 61.070 104.800 ;
        RECT 61.250 104.750 62.250 105.085 ;
        RECT 82.305 104.800 82.495 105.345 ;
        RECT 83.905 105.240 84.095 105.345 ;
        RECT 86.570 105.340 86.800 106.860 ;
        RECT 87.160 105.340 87.390 106.860 ;
        RECT 83.905 105.085 84.910 105.240 ;
        RECT 86.570 105.150 87.390 105.340 ;
        RECT 86.570 105.100 86.800 105.150 ;
        RECT 87.160 105.100 87.390 105.150 ;
        RECT 92.800 105.100 93.030 106.860 ;
        RECT 94.680 105.100 94.910 106.860 ;
        RECT 96.465 106.855 96.790 107.100 ;
        RECT 96.560 105.100 96.790 106.855 ;
        RECT 98.325 107.055 98.515 108.150 ;
        RECT 99.280 108.060 99.550 108.150 ;
        RECT 99.320 107.155 99.510 107.185 ;
        RECT 99.280 107.055 99.550 107.155 ;
        RECT 109.350 107.100 109.915 108.190 ;
        RECT 115.375 107.100 115.565 108.190 ;
        RECT 117.245 107.100 117.435 108.190 ;
        RECT 119.125 107.100 119.315 108.190 ;
        RECT 120.985 108.150 122.210 108.340 ;
        RECT 98.325 106.865 99.550 107.055 ;
        RECT 98.325 105.770 98.515 106.865 ;
        RECT 99.280 106.775 99.550 106.865 ;
        RECT 109.230 106.860 110.050 107.100 ;
        RECT 115.375 106.860 115.690 107.100 ;
        RECT 117.245 106.860 117.570 107.100 ;
        RECT 99.320 105.870 99.510 105.905 ;
        RECT 99.280 105.770 99.550 105.870 ;
        RECT 98.325 105.580 99.550 105.770 ;
        RECT 99.280 105.490 99.550 105.580 ;
        RECT 103.770 105.405 106.755 105.535 ;
        RECT 103.415 105.345 106.755 105.405 ;
        RECT 103.415 105.195 103.970 105.345 ;
        RECT 103.415 105.175 103.705 105.195 ;
        RECT 59.440 104.300 59.670 104.610 ;
        RECT 60.840 104.560 62.250 104.750 ;
        RECT 60.840 104.300 61.070 104.560 ;
        RECT 61.250 104.240 62.250 104.560 ;
        RECT 82.100 104.610 82.495 104.800 ;
        RECT 83.500 104.750 83.730 104.800 ;
        RECT 83.910 104.750 84.910 105.085 ;
        RECT 104.965 104.800 105.155 105.345 ;
        RECT 106.565 105.240 106.755 105.345 ;
        RECT 109.230 105.340 109.460 106.860 ;
        RECT 109.820 105.340 110.050 106.860 ;
        RECT 106.565 105.085 107.570 105.240 ;
        RECT 109.230 105.150 110.050 105.340 ;
        RECT 109.230 105.100 109.460 105.150 ;
        RECT 109.820 105.100 110.050 105.150 ;
        RECT 115.460 105.100 115.690 106.860 ;
        RECT 117.340 105.100 117.570 106.860 ;
        RECT 119.125 106.855 119.450 107.100 ;
        RECT 119.220 105.100 119.450 106.855 ;
        RECT 120.985 107.055 121.175 108.150 ;
        RECT 121.940 108.060 122.210 108.150 ;
        RECT 121.980 107.155 122.170 107.185 ;
        RECT 121.940 107.055 122.210 107.155 ;
        RECT 120.985 106.865 122.210 107.055 ;
        RECT 120.985 105.770 121.175 106.865 ;
        RECT 121.940 106.775 122.210 106.865 ;
        RECT 121.980 105.870 122.170 105.905 ;
        RECT 121.940 105.770 122.210 105.870 ;
        RECT 120.985 105.580 122.210 105.770 ;
        RECT 121.940 105.490 122.210 105.580 ;
        RECT 82.100 104.300 82.330 104.610 ;
        RECT 83.500 104.560 84.910 104.750 ;
        RECT 83.500 104.300 83.730 104.560 ;
        RECT 83.910 104.240 84.910 104.560 ;
        RECT 104.760 104.610 105.155 104.800 ;
        RECT 106.160 104.750 106.390 104.800 ;
        RECT 106.570 104.750 107.570 105.085 ;
        RECT 104.760 104.300 104.990 104.610 ;
        RECT 106.160 104.560 107.570 104.750 ;
        RECT 106.160 104.300 106.390 104.560 ;
        RECT 106.570 104.240 107.570 104.560 ;
        RECT 41.250 92.820 41.480 92.850 ;
        RECT 41.840 92.820 42.070 92.850 ;
        RECT 41.250 92.220 42.070 92.820 ;
        RECT 47.400 92.250 48.000 92.850 ;
        RECT 49.280 92.250 49.880 92.850 ;
        RECT 51.160 92.250 51.760 92.850 ;
        RECT 63.910 92.820 64.140 92.850 ;
        RECT 64.500 92.820 64.730 92.850 ;
        RECT 52.970 92.340 53.230 92.660 ;
        RECT 54.000 92.390 54.190 92.420 ;
        RECT 53.005 92.290 53.230 92.340 ;
        RECT 53.960 92.290 54.230 92.390 ;
        RECT 41.250 91.100 41.480 92.220 ;
        RECT 41.840 91.100 42.070 92.220 ;
        RECT 41.250 90.850 42.070 91.100 ;
        RECT 47.480 91.095 47.710 92.250 ;
        RECT 49.360 91.105 49.590 92.250 ;
        RECT 51.240 91.105 51.470 92.250 ;
        RECT 47.395 90.850 47.710 91.095 ;
        RECT 49.265 90.850 49.590 91.105 ;
        RECT 51.145 90.850 51.470 91.105 ;
        RECT 53.005 92.100 54.230 92.290 ;
        RECT 53.005 91.000 53.195 92.100 ;
        RECT 53.960 92.010 54.230 92.100 ;
        RECT 63.910 92.220 64.730 92.820 ;
        RECT 70.060 92.250 70.660 92.850 ;
        RECT 71.940 92.250 72.540 92.850 ;
        RECT 73.820 92.250 74.420 92.850 ;
        RECT 86.570 92.820 86.800 92.850 ;
        RECT 87.160 92.820 87.390 92.850 ;
        RECT 75.630 92.340 75.890 92.660 ;
        RECT 76.660 92.390 76.850 92.420 ;
        RECT 75.665 92.290 75.890 92.340 ;
        RECT 76.620 92.290 76.890 92.390 ;
        RECT 54.000 91.100 54.190 91.130 ;
        RECT 63.910 91.100 64.140 92.220 ;
        RECT 64.500 91.100 64.730 92.220 ;
        RECT 53.960 91.000 54.230 91.100 ;
        RECT 41.370 89.760 41.935 90.850 ;
        RECT 47.395 89.760 47.585 90.850 ;
        RECT 49.265 89.760 49.455 90.850 ;
        RECT 51.145 89.760 51.335 90.850 ;
        RECT 53.005 90.810 54.230 91.000 ;
        RECT 63.910 90.850 64.730 91.100 ;
        RECT 70.140 91.095 70.370 92.250 ;
        RECT 72.020 91.105 72.250 92.250 ;
        RECT 73.900 91.105 74.130 92.250 ;
        RECT 70.055 90.850 70.370 91.095 ;
        RECT 71.925 90.850 72.250 91.105 ;
        RECT 73.805 90.850 74.130 91.105 ;
        RECT 75.665 92.100 76.890 92.290 ;
        RECT 75.665 91.000 75.855 92.100 ;
        RECT 76.620 92.010 76.890 92.100 ;
        RECT 86.570 92.220 87.390 92.820 ;
        RECT 92.720 92.250 93.320 92.850 ;
        RECT 94.600 92.250 95.200 92.850 ;
        RECT 96.480 92.250 97.080 92.850 ;
        RECT 109.230 92.820 109.460 92.850 ;
        RECT 109.820 92.820 110.050 92.850 ;
        RECT 98.290 92.340 98.550 92.660 ;
        RECT 99.320 92.390 99.510 92.420 ;
        RECT 98.325 92.290 98.550 92.340 ;
        RECT 99.280 92.290 99.550 92.390 ;
        RECT 76.660 91.100 76.850 91.130 ;
        RECT 86.570 91.100 86.800 92.220 ;
        RECT 87.160 91.100 87.390 92.220 ;
        RECT 76.620 91.000 76.890 91.100 ;
        RECT 41.250 89.520 42.070 89.760 ;
        RECT 47.395 89.520 47.710 89.760 ;
        RECT 49.265 89.520 49.590 89.760 ;
        RECT 35.790 88.065 38.775 88.195 ;
        RECT 35.435 88.005 38.775 88.065 ;
        RECT 35.435 87.855 35.990 88.005 ;
        RECT 35.435 87.835 35.725 87.855 ;
        RECT 36.985 87.460 37.175 88.005 ;
        RECT 38.585 87.900 38.775 88.005 ;
        RECT 41.250 88.000 41.480 89.520 ;
        RECT 41.840 88.000 42.070 89.520 ;
        RECT 38.585 87.745 39.590 87.900 ;
        RECT 41.250 87.810 42.070 88.000 ;
        RECT 41.250 87.760 41.480 87.810 ;
        RECT 41.840 87.760 42.070 87.810 ;
        RECT 47.480 87.760 47.710 89.520 ;
        RECT 49.360 87.760 49.590 89.520 ;
        RECT 51.145 89.515 51.470 89.760 ;
        RECT 51.240 87.760 51.470 89.515 ;
        RECT 53.005 89.715 53.195 90.810 ;
        RECT 53.960 90.720 54.230 90.810 ;
        RECT 54.000 89.815 54.190 89.845 ;
        RECT 53.960 89.715 54.230 89.815 ;
        RECT 64.030 89.760 64.595 90.850 ;
        RECT 70.055 89.760 70.245 90.850 ;
        RECT 71.925 89.760 72.115 90.850 ;
        RECT 73.805 89.760 73.995 90.850 ;
        RECT 75.665 90.810 76.890 91.000 ;
        RECT 86.570 90.850 87.390 91.100 ;
        RECT 92.800 91.095 93.030 92.250 ;
        RECT 94.680 91.105 94.910 92.250 ;
        RECT 96.560 91.105 96.790 92.250 ;
        RECT 92.715 90.850 93.030 91.095 ;
        RECT 94.585 90.850 94.910 91.105 ;
        RECT 96.465 90.850 96.790 91.105 ;
        RECT 98.325 92.100 99.550 92.290 ;
        RECT 98.325 91.000 98.515 92.100 ;
        RECT 99.280 92.010 99.550 92.100 ;
        RECT 109.230 92.220 110.050 92.820 ;
        RECT 115.380 92.250 115.980 92.850 ;
        RECT 117.260 92.250 117.860 92.850 ;
        RECT 119.140 92.250 119.740 92.850 ;
        RECT 120.950 92.340 121.210 92.660 ;
        RECT 121.980 92.390 122.170 92.420 ;
        RECT 120.985 92.290 121.210 92.340 ;
        RECT 121.940 92.290 122.210 92.390 ;
        RECT 99.320 91.100 99.510 91.130 ;
        RECT 109.230 91.100 109.460 92.220 ;
        RECT 109.820 91.100 110.050 92.220 ;
        RECT 99.280 91.000 99.550 91.100 ;
        RECT 53.005 89.525 54.230 89.715 ;
        RECT 53.005 88.430 53.195 89.525 ;
        RECT 53.960 89.435 54.230 89.525 ;
        RECT 63.910 89.520 64.730 89.760 ;
        RECT 70.055 89.520 70.370 89.760 ;
        RECT 71.925 89.520 72.250 89.760 ;
        RECT 54.000 88.530 54.190 88.565 ;
        RECT 53.960 88.430 54.230 88.530 ;
        RECT 53.005 88.240 54.230 88.430 ;
        RECT 53.960 88.150 54.230 88.240 ;
        RECT 58.450 88.065 61.435 88.195 ;
        RECT 58.095 88.005 61.435 88.065 ;
        RECT 58.095 87.855 58.650 88.005 ;
        RECT 58.095 87.835 58.385 87.855 ;
        RECT 36.780 87.270 37.175 87.460 ;
        RECT 38.180 87.410 38.410 87.460 ;
        RECT 38.590 87.410 39.590 87.745 ;
        RECT 59.645 87.460 59.835 88.005 ;
        RECT 61.245 87.900 61.435 88.005 ;
        RECT 63.910 88.000 64.140 89.520 ;
        RECT 64.500 88.000 64.730 89.520 ;
        RECT 61.245 87.745 62.250 87.900 ;
        RECT 63.910 87.810 64.730 88.000 ;
        RECT 63.910 87.760 64.140 87.810 ;
        RECT 64.500 87.760 64.730 87.810 ;
        RECT 70.140 87.760 70.370 89.520 ;
        RECT 72.020 87.760 72.250 89.520 ;
        RECT 73.805 89.515 74.130 89.760 ;
        RECT 73.900 87.760 74.130 89.515 ;
        RECT 75.665 89.715 75.855 90.810 ;
        RECT 76.620 90.720 76.890 90.810 ;
        RECT 76.660 89.815 76.850 89.845 ;
        RECT 76.620 89.715 76.890 89.815 ;
        RECT 86.690 89.760 87.255 90.850 ;
        RECT 92.715 89.760 92.905 90.850 ;
        RECT 94.585 89.760 94.775 90.850 ;
        RECT 96.465 89.760 96.655 90.850 ;
        RECT 98.325 90.810 99.550 91.000 ;
        RECT 109.230 90.850 110.050 91.100 ;
        RECT 115.460 91.095 115.690 92.250 ;
        RECT 117.340 91.105 117.570 92.250 ;
        RECT 119.220 91.105 119.450 92.250 ;
        RECT 115.375 90.850 115.690 91.095 ;
        RECT 117.245 90.850 117.570 91.105 ;
        RECT 119.125 90.850 119.450 91.105 ;
        RECT 120.985 92.100 122.210 92.290 ;
        RECT 120.985 91.000 121.175 92.100 ;
        RECT 121.940 92.010 122.210 92.100 ;
        RECT 121.980 91.100 122.170 91.130 ;
        RECT 121.940 91.000 122.210 91.100 ;
        RECT 75.665 89.525 76.890 89.715 ;
        RECT 75.665 88.430 75.855 89.525 ;
        RECT 76.620 89.435 76.890 89.525 ;
        RECT 86.570 89.520 87.390 89.760 ;
        RECT 92.715 89.520 93.030 89.760 ;
        RECT 94.585 89.520 94.910 89.760 ;
        RECT 76.660 88.530 76.850 88.565 ;
        RECT 76.620 88.430 76.890 88.530 ;
        RECT 75.665 88.240 76.890 88.430 ;
        RECT 76.620 88.150 76.890 88.240 ;
        RECT 81.110 88.065 84.095 88.195 ;
        RECT 80.755 88.005 84.095 88.065 ;
        RECT 80.755 87.855 81.310 88.005 ;
        RECT 80.755 87.835 81.045 87.855 ;
        RECT 36.780 86.960 37.010 87.270 ;
        RECT 38.180 87.220 39.590 87.410 ;
        RECT 38.180 86.960 38.410 87.220 ;
        RECT 38.590 86.900 39.590 87.220 ;
        RECT 59.440 87.270 59.835 87.460 ;
        RECT 60.840 87.410 61.070 87.460 ;
        RECT 61.250 87.410 62.250 87.745 ;
        RECT 82.305 87.460 82.495 88.005 ;
        RECT 83.905 87.900 84.095 88.005 ;
        RECT 86.570 88.000 86.800 89.520 ;
        RECT 87.160 88.000 87.390 89.520 ;
        RECT 83.905 87.745 84.910 87.900 ;
        RECT 86.570 87.810 87.390 88.000 ;
        RECT 86.570 87.760 86.800 87.810 ;
        RECT 87.160 87.760 87.390 87.810 ;
        RECT 92.800 87.760 93.030 89.520 ;
        RECT 94.680 87.760 94.910 89.520 ;
        RECT 96.465 89.515 96.790 89.760 ;
        RECT 96.560 87.760 96.790 89.515 ;
        RECT 98.325 89.715 98.515 90.810 ;
        RECT 99.280 90.720 99.550 90.810 ;
        RECT 99.320 89.815 99.510 89.845 ;
        RECT 99.280 89.715 99.550 89.815 ;
        RECT 109.350 89.760 109.915 90.850 ;
        RECT 115.375 89.760 115.565 90.850 ;
        RECT 117.245 89.760 117.435 90.850 ;
        RECT 119.125 89.760 119.315 90.850 ;
        RECT 120.985 90.810 122.210 91.000 ;
        RECT 98.325 89.525 99.550 89.715 ;
        RECT 98.325 88.430 98.515 89.525 ;
        RECT 99.280 89.435 99.550 89.525 ;
        RECT 109.230 89.520 110.050 89.760 ;
        RECT 115.375 89.520 115.690 89.760 ;
        RECT 117.245 89.520 117.570 89.760 ;
        RECT 99.320 88.530 99.510 88.565 ;
        RECT 99.280 88.430 99.550 88.530 ;
        RECT 98.325 88.240 99.550 88.430 ;
        RECT 99.280 88.150 99.550 88.240 ;
        RECT 103.770 88.065 106.755 88.195 ;
        RECT 103.415 88.005 106.755 88.065 ;
        RECT 103.415 87.855 103.970 88.005 ;
        RECT 103.415 87.835 103.705 87.855 ;
        RECT 59.440 86.960 59.670 87.270 ;
        RECT 60.840 87.220 62.250 87.410 ;
        RECT 60.840 86.960 61.070 87.220 ;
        RECT 61.250 86.900 62.250 87.220 ;
        RECT 82.100 87.270 82.495 87.460 ;
        RECT 83.500 87.410 83.730 87.460 ;
        RECT 83.910 87.410 84.910 87.745 ;
        RECT 104.965 87.460 105.155 88.005 ;
        RECT 106.565 87.900 106.755 88.005 ;
        RECT 109.230 88.000 109.460 89.520 ;
        RECT 109.820 88.000 110.050 89.520 ;
        RECT 106.565 87.745 107.570 87.900 ;
        RECT 109.230 87.810 110.050 88.000 ;
        RECT 109.230 87.760 109.460 87.810 ;
        RECT 109.820 87.760 110.050 87.810 ;
        RECT 115.460 87.760 115.690 89.520 ;
        RECT 117.340 87.760 117.570 89.520 ;
        RECT 119.125 89.515 119.450 89.760 ;
        RECT 119.220 87.760 119.450 89.515 ;
        RECT 120.985 89.715 121.175 90.810 ;
        RECT 121.940 90.720 122.210 90.810 ;
        RECT 121.980 89.815 122.170 89.845 ;
        RECT 121.940 89.715 122.210 89.815 ;
        RECT 120.985 89.525 122.210 89.715 ;
        RECT 120.985 88.430 121.175 89.525 ;
        RECT 121.940 89.435 122.210 89.525 ;
        RECT 121.980 88.530 122.170 88.565 ;
        RECT 121.940 88.430 122.210 88.530 ;
        RECT 120.985 88.240 122.210 88.430 ;
        RECT 121.940 88.150 122.210 88.240 ;
        RECT 82.100 86.960 82.330 87.270 ;
        RECT 83.500 87.220 84.910 87.410 ;
        RECT 83.500 86.960 83.730 87.220 ;
        RECT 83.910 86.900 84.910 87.220 ;
        RECT 104.760 87.270 105.155 87.460 ;
        RECT 106.160 87.410 106.390 87.460 ;
        RECT 106.570 87.410 107.570 87.745 ;
        RECT 104.760 86.960 104.990 87.270 ;
        RECT 106.160 87.220 107.570 87.410 ;
        RECT 106.160 86.960 106.390 87.220 ;
        RECT 106.570 86.900 107.570 87.220 ;
        RECT 41.250 75.480 41.480 75.510 ;
        RECT 41.840 75.480 42.070 75.510 ;
        RECT 41.250 74.880 42.070 75.480 ;
        RECT 47.400 74.910 48.000 75.510 ;
        RECT 49.280 74.910 49.880 75.510 ;
        RECT 51.160 74.910 51.760 75.510 ;
        RECT 63.910 75.480 64.140 75.510 ;
        RECT 64.500 75.480 64.730 75.510 ;
        RECT 52.970 75.000 53.230 75.320 ;
        RECT 54.000 75.050 54.190 75.080 ;
        RECT 53.005 74.950 53.230 75.000 ;
        RECT 53.960 74.950 54.230 75.050 ;
        RECT 41.250 73.760 41.480 74.880 ;
        RECT 41.840 73.760 42.070 74.880 ;
        RECT 41.250 73.510 42.070 73.760 ;
        RECT 47.480 73.755 47.710 74.910 ;
        RECT 49.360 73.765 49.590 74.910 ;
        RECT 51.240 73.765 51.470 74.910 ;
        RECT 47.395 73.510 47.710 73.755 ;
        RECT 49.265 73.510 49.590 73.765 ;
        RECT 51.145 73.510 51.470 73.765 ;
        RECT 53.005 74.760 54.230 74.950 ;
        RECT 53.005 73.660 53.195 74.760 ;
        RECT 53.960 74.670 54.230 74.760 ;
        RECT 63.910 74.880 64.730 75.480 ;
        RECT 70.060 74.910 70.660 75.510 ;
        RECT 71.940 74.910 72.540 75.510 ;
        RECT 73.820 74.910 74.420 75.510 ;
        RECT 86.570 75.480 86.800 75.510 ;
        RECT 87.160 75.480 87.390 75.510 ;
        RECT 75.630 75.000 75.890 75.320 ;
        RECT 76.660 75.050 76.850 75.080 ;
        RECT 75.665 74.950 75.890 75.000 ;
        RECT 76.620 74.950 76.890 75.050 ;
        RECT 54.000 73.760 54.190 73.790 ;
        RECT 63.910 73.760 64.140 74.880 ;
        RECT 64.500 73.760 64.730 74.880 ;
        RECT 53.960 73.660 54.230 73.760 ;
        RECT 41.370 72.420 41.935 73.510 ;
        RECT 47.395 72.420 47.585 73.510 ;
        RECT 49.265 72.420 49.455 73.510 ;
        RECT 51.145 72.420 51.335 73.510 ;
        RECT 53.005 73.470 54.230 73.660 ;
        RECT 63.910 73.510 64.730 73.760 ;
        RECT 70.140 73.755 70.370 74.910 ;
        RECT 72.020 73.765 72.250 74.910 ;
        RECT 73.900 73.765 74.130 74.910 ;
        RECT 70.055 73.510 70.370 73.755 ;
        RECT 71.925 73.510 72.250 73.765 ;
        RECT 73.805 73.510 74.130 73.765 ;
        RECT 75.665 74.760 76.890 74.950 ;
        RECT 75.665 73.660 75.855 74.760 ;
        RECT 76.620 74.670 76.890 74.760 ;
        RECT 86.570 74.880 87.390 75.480 ;
        RECT 92.720 74.910 93.320 75.510 ;
        RECT 94.600 74.910 95.200 75.510 ;
        RECT 96.480 74.910 97.080 75.510 ;
        RECT 109.230 75.480 109.460 75.510 ;
        RECT 109.820 75.480 110.050 75.510 ;
        RECT 98.290 75.000 98.550 75.320 ;
        RECT 99.320 75.050 99.510 75.080 ;
        RECT 98.325 74.950 98.550 75.000 ;
        RECT 99.280 74.950 99.550 75.050 ;
        RECT 76.660 73.760 76.850 73.790 ;
        RECT 86.570 73.760 86.800 74.880 ;
        RECT 87.160 73.760 87.390 74.880 ;
        RECT 76.620 73.660 76.890 73.760 ;
        RECT 41.250 72.180 42.070 72.420 ;
        RECT 47.395 72.180 47.710 72.420 ;
        RECT 49.265 72.180 49.590 72.420 ;
        RECT 35.790 70.725 38.775 70.855 ;
        RECT 35.435 70.665 38.775 70.725 ;
        RECT 35.435 70.515 35.990 70.665 ;
        RECT 35.435 70.495 35.725 70.515 ;
        RECT 36.985 70.120 37.175 70.665 ;
        RECT 38.585 70.560 38.775 70.665 ;
        RECT 41.250 70.660 41.480 72.180 ;
        RECT 41.840 70.660 42.070 72.180 ;
        RECT 38.585 70.405 39.590 70.560 ;
        RECT 41.250 70.470 42.070 70.660 ;
        RECT 41.250 70.420 41.480 70.470 ;
        RECT 41.840 70.420 42.070 70.470 ;
        RECT 47.480 70.420 47.710 72.180 ;
        RECT 49.360 70.420 49.590 72.180 ;
        RECT 51.145 72.175 51.470 72.420 ;
        RECT 51.240 70.420 51.470 72.175 ;
        RECT 53.005 72.375 53.195 73.470 ;
        RECT 53.960 73.380 54.230 73.470 ;
        RECT 54.000 72.475 54.190 72.505 ;
        RECT 53.960 72.375 54.230 72.475 ;
        RECT 64.030 72.420 64.595 73.510 ;
        RECT 70.055 72.420 70.245 73.510 ;
        RECT 71.925 72.420 72.115 73.510 ;
        RECT 73.805 72.420 73.995 73.510 ;
        RECT 75.665 73.470 76.890 73.660 ;
        RECT 86.570 73.510 87.390 73.760 ;
        RECT 92.800 73.755 93.030 74.910 ;
        RECT 94.680 73.765 94.910 74.910 ;
        RECT 96.560 73.765 96.790 74.910 ;
        RECT 92.715 73.510 93.030 73.755 ;
        RECT 94.585 73.510 94.910 73.765 ;
        RECT 96.465 73.510 96.790 73.765 ;
        RECT 98.325 74.760 99.550 74.950 ;
        RECT 98.325 73.660 98.515 74.760 ;
        RECT 99.280 74.670 99.550 74.760 ;
        RECT 109.230 74.880 110.050 75.480 ;
        RECT 115.380 74.910 115.980 75.510 ;
        RECT 117.260 74.910 117.860 75.510 ;
        RECT 119.140 74.910 119.740 75.510 ;
        RECT 120.950 75.000 121.210 75.320 ;
        RECT 121.980 75.050 122.170 75.080 ;
        RECT 120.985 74.950 121.210 75.000 ;
        RECT 121.940 74.950 122.210 75.050 ;
        RECT 99.320 73.760 99.510 73.790 ;
        RECT 109.230 73.760 109.460 74.880 ;
        RECT 109.820 73.760 110.050 74.880 ;
        RECT 99.280 73.660 99.550 73.760 ;
        RECT 53.005 72.185 54.230 72.375 ;
        RECT 53.005 71.090 53.195 72.185 ;
        RECT 53.960 72.095 54.230 72.185 ;
        RECT 63.910 72.180 64.730 72.420 ;
        RECT 70.055 72.180 70.370 72.420 ;
        RECT 71.925 72.180 72.250 72.420 ;
        RECT 54.000 71.190 54.190 71.225 ;
        RECT 53.960 71.090 54.230 71.190 ;
        RECT 53.005 70.900 54.230 71.090 ;
        RECT 53.960 70.810 54.230 70.900 ;
        RECT 58.450 70.725 61.435 70.855 ;
        RECT 58.095 70.665 61.435 70.725 ;
        RECT 58.095 70.515 58.650 70.665 ;
        RECT 58.095 70.495 58.385 70.515 ;
        RECT 36.780 69.930 37.175 70.120 ;
        RECT 38.180 70.070 38.410 70.120 ;
        RECT 38.590 70.070 39.590 70.405 ;
        RECT 59.645 70.120 59.835 70.665 ;
        RECT 61.245 70.560 61.435 70.665 ;
        RECT 63.910 70.660 64.140 72.180 ;
        RECT 64.500 70.660 64.730 72.180 ;
        RECT 61.245 70.405 62.250 70.560 ;
        RECT 63.910 70.470 64.730 70.660 ;
        RECT 63.910 70.420 64.140 70.470 ;
        RECT 64.500 70.420 64.730 70.470 ;
        RECT 70.140 70.420 70.370 72.180 ;
        RECT 72.020 70.420 72.250 72.180 ;
        RECT 73.805 72.175 74.130 72.420 ;
        RECT 73.900 70.420 74.130 72.175 ;
        RECT 75.665 72.375 75.855 73.470 ;
        RECT 76.620 73.380 76.890 73.470 ;
        RECT 76.660 72.475 76.850 72.505 ;
        RECT 76.620 72.375 76.890 72.475 ;
        RECT 86.690 72.420 87.255 73.510 ;
        RECT 92.715 72.420 92.905 73.510 ;
        RECT 94.585 72.420 94.775 73.510 ;
        RECT 96.465 72.420 96.655 73.510 ;
        RECT 98.325 73.470 99.550 73.660 ;
        RECT 109.230 73.510 110.050 73.760 ;
        RECT 115.460 73.755 115.690 74.910 ;
        RECT 117.340 73.765 117.570 74.910 ;
        RECT 119.220 73.765 119.450 74.910 ;
        RECT 115.375 73.510 115.690 73.755 ;
        RECT 117.245 73.510 117.570 73.765 ;
        RECT 119.125 73.510 119.450 73.765 ;
        RECT 120.985 74.760 122.210 74.950 ;
        RECT 120.985 73.660 121.175 74.760 ;
        RECT 121.940 74.670 122.210 74.760 ;
        RECT 121.980 73.760 122.170 73.790 ;
        RECT 121.940 73.660 122.210 73.760 ;
        RECT 75.665 72.185 76.890 72.375 ;
        RECT 75.665 71.090 75.855 72.185 ;
        RECT 76.620 72.095 76.890 72.185 ;
        RECT 86.570 72.180 87.390 72.420 ;
        RECT 92.715 72.180 93.030 72.420 ;
        RECT 94.585 72.180 94.910 72.420 ;
        RECT 76.660 71.190 76.850 71.225 ;
        RECT 76.620 71.090 76.890 71.190 ;
        RECT 75.665 70.900 76.890 71.090 ;
        RECT 76.620 70.810 76.890 70.900 ;
        RECT 81.110 70.725 84.095 70.855 ;
        RECT 80.755 70.665 84.095 70.725 ;
        RECT 80.755 70.515 81.310 70.665 ;
        RECT 80.755 70.495 81.045 70.515 ;
        RECT 36.780 69.620 37.010 69.930 ;
        RECT 38.180 69.880 39.590 70.070 ;
        RECT 38.180 69.620 38.410 69.880 ;
        RECT 38.590 69.560 39.590 69.880 ;
        RECT 59.440 69.930 59.835 70.120 ;
        RECT 60.840 70.070 61.070 70.120 ;
        RECT 61.250 70.070 62.250 70.405 ;
        RECT 82.305 70.120 82.495 70.665 ;
        RECT 83.905 70.560 84.095 70.665 ;
        RECT 86.570 70.660 86.800 72.180 ;
        RECT 87.160 70.660 87.390 72.180 ;
        RECT 83.905 70.405 84.910 70.560 ;
        RECT 86.570 70.470 87.390 70.660 ;
        RECT 86.570 70.420 86.800 70.470 ;
        RECT 87.160 70.420 87.390 70.470 ;
        RECT 92.800 70.420 93.030 72.180 ;
        RECT 94.680 70.420 94.910 72.180 ;
        RECT 96.465 72.175 96.790 72.420 ;
        RECT 96.560 70.420 96.790 72.175 ;
        RECT 98.325 72.375 98.515 73.470 ;
        RECT 99.280 73.380 99.550 73.470 ;
        RECT 99.320 72.475 99.510 72.505 ;
        RECT 99.280 72.375 99.550 72.475 ;
        RECT 109.350 72.420 109.915 73.510 ;
        RECT 115.375 72.420 115.565 73.510 ;
        RECT 117.245 72.420 117.435 73.510 ;
        RECT 119.125 72.420 119.315 73.510 ;
        RECT 120.985 73.470 122.210 73.660 ;
        RECT 98.325 72.185 99.550 72.375 ;
        RECT 98.325 71.090 98.515 72.185 ;
        RECT 99.280 72.095 99.550 72.185 ;
        RECT 109.230 72.180 110.050 72.420 ;
        RECT 115.375 72.180 115.690 72.420 ;
        RECT 117.245 72.180 117.570 72.420 ;
        RECT 99.320 71.190 99.510 71.225 ;
        RECT 99.280 71.090 99.550 71.190 ;
        RECT 98.325 70.900 99.550 71.090 ;
        RECT 99.280 70.810 99.550 70.900 ;
        RECT 103.770 70.725 106.755 70.855 ;
        RECT 103.415 70.665 106.755 70.725 ;
        RECT 103.415 70.515 103.970 70.665 ;
        RECT 103.415 70.495 103.705 70.515 ;
        RECT 59.440 69.620 59.670 69.930 ;
        RECT 60.840 69.880 62.250 70.070 ;
        RECT 60.840 69.620 61.070 69.880 ;
        RECT 61.250 69.560 62.250 69.880 ;
        RECT 82.100 69.930 82.495 70.120 ;
        RECT 83.500 70.070 83.730 70.120 ;
        RECT 83.910 70.070 84.910 70.405 ;
        RECT 104.965 70.120 105.155 70.665 ;
        RECT 106.565 70.560 106.755 70.665 ;
        RECT 109.230 70.660 109.460 72.180 ;
        RECT 109.820 70.660 110.050 72.180 ;
        RECT 106.565 70.405 107.570 70.560 ;
        RECT 109.230 70.470 110.050 70.660 ;
        RECT 109.230 70.420 109.460 70.470 ;
        RECT 109.820 70.420 110.050 70.470 ;
        RECT 115.460 70.420 115.690 72.180 ;
        RECT 117.340 70.420 117.570 72.180 ;
        RECT 119.125 72.175 119.450 72.420 ;
        RECT 119.220 70.420 119.450 72.175 ;
        RECT 120.985 72.375 121.175 73.470 ;
        RECT 121.940 73.380 122.210 73.470 ;
        RECT 121.980 72.475 122.170 72.505 ;
        RECT 121.940 72.375 122.210 72.475 ;
        RECT 120.985 72.185 122.210 72.375 ;
        RECT 120.985 71.090 121.175 72.185 ;
        RECT 121.940 72.095 122.210 72.185 ;
        RECT 121.980 71.190 122.170 71.225 ;
        RECT 121.940 71.090 122.210 71.190 ;
        RECT 120.985 70.900 122.210 71.090 ;
        RECT 121.940 70.810 122.210 70.900 ;
        RECT 82.100 69.620 82.330 69.930 ;
        RECT 83.500 69.880 84.910 70.070 ;
        RECT 83.500 69.620 83.730 69.880 ;
        RECT 83.910 69.560 84.910 69.880 ;
        RECT 104.760 69.930 105.155 70.120 ;
        RECT 106.160 70.070 106.390 70.120 ;
        RECT 106.570 70.070 107.570 70.405 ;
        RECT 104.760 69.620 104.990 69.930 ;
        RECT 106.160 69.880 107.570 70.070 ;
        RECT 106.160 69.620 106.390 69.880 ;
        RECT 106.570 69.560 107.570 69.880 ;
        RECT 41.250 57.480 41.480 57.510 ;
        RECT 41.840 57.480 42.070 57.510 ;
        RECT 41.250 56.880 42.070 57.480 ;
        RECT 47.400 56.910 48.000 57.510 ;
        RECT 49.280 56.910 49.880 57.510 ;
        RECT 51.160 56.910 51.760 57.510 ;
        RECT 63.910 57.480 64.140 57.510 ;
        RECT 64.500 57.480 64.730 57.510 ;
        RECT 52.970 57.000 53.230 57.320 ;
        RECT 54.000 57.050 54.190 57.080 ;
        RECT 53.005 56.950 53.230 57.000 ;
        RECT 53.960 56.950 54.230 57.050 ;
        RECT 41.250 55.760 41.480 56.880 ;
        RECT 41.840 55.760 42.070 56.880 ;
        RECT 41.250 55.510 42.070 55.760 ;
        RECT 47.480 55.755 47.710 56.910 ;
        RECT 49.360 55.765 49.590 56.910 ;
        RECT 51.240 55.765 51.470 56.910 ;
        RECT 47.395 55.510 47.710 55.755 ;
        RECT 49.265 55.510 49.590 55.765 ;
        RECT 51.145 55.510 51.470 55.765 ;
        RECT 53.005 56.760 54.230 56.950 ;
        RECT 53.005 55.660 53.195 56.760 ;
        RECT 53.960 56.670 54.230 56.760 ;
        RECT 63.910 56.880 64.730 57.480 ;
        RECT 70.060 56.910 70.660 57.510 ;
        RECT 71.940 56.910 72.540 57.510 ;
        RECT 73.820 56.910 74.420 57.510 ;
        RECT 86.570 57.480 86.800 57.510 ;
        RECT 87.160 57.480 87.390 57.510 ;
        RECT 75.630 57.000 75.890 57.320 ;
        RECT 76.660 57.050 76.850 57.080 ;
        RECT 75.665 56.950 75.890 57.000 ;
        RECT 76.620 56.950 76.890 57.050 ;
        RECT 54.000 55.760 54.190 55.790 ;
        RECT 63.910 55.760 64.140 56.880 ;
        RECT 64.500 55.760 64.730 56.880 ;
        RECT 53.960 55.660 54.230 55.760 ;
        RECT 41.370 54.420 41.935 55.510 ;
        RECT 47.395 54.420 47.585 55.510 ;
        RECT 49.265 54.420 49.455 55.510 ;
        RECT 51.145 54.420 51.335 55.510 ;
        RECT 53.005 55.470 54.230 55.660 ;
        RECT 63.910 55.510 64.730 55.760 ;
        RECT 70.140 55.755 70.370 56.910 ;
        RECT 72.020 55.765 72.250 56.910 ;
        RECT 73.900 55.765 74.130 56.910 ;
        RECT 70.055 55.510 70.370 55.755 ;
        RECT 71.925 55.510 72.250 55.765 ;
        RECT 73.805 55.510 74.130 55.765 ;
        RECT 75.665 56.760 76.890 56.950 ;
        RECT 75.665 55.660 75.855 56.760 ;
        RECT 76.620 56.670 76.890 56.760 ;
        RECT 86.570 56.880 87.390 57.480 ;
        RECT 92.720 56.910 93.320 57.510 ;
        RECT 94.600 56.910 95.200 57.510 ;
        RECT 96.480 56.910 97.080 57.510 ;
        RECT 109.230 57.480 109.460 57.510 ;
        RECT 109.820 57.480 110.050 57.510 ;
        RECT 98.290 57.000 98.550 57.320 ;
        RECT 99.320 57.050 99.510 57.080 ;
        RECT 98.325 56.950 98.550 57.000 ;
        RECT 99.280 56.950 99.550 57.050 ;
        RECT 76.660 55.760 76.850 55.790 ;
        RECT 86.570 55.760 86.800 56.880 ;
        RECT 87.160 55.760 87.390 56.880 ;
        RECT 76.620 55.660 76.890 55.760 ;
        RECT 41.250 54.180 42.070 54.420 ;
        RECT 47.395 54.180 47.710 54.420 ;
        RECT 49.265 54.180 49.590 54.420 ;
        RECT 41.250 52.660 41.480 54.180 ;
        RECT 41.840 52.660 42.070 54.180 ;
        RECT 41.250 52.470 42.070 52.660 ;
        RECT 41.250 52.420 41.480 52.470 ;
        RECT 41.840 52.420 42.070 52.470 ;
        RECT 47.480 52.420 47.710 54.180 ;
        RECT 49.360 52.420 49.590 54.180 ;
        RECT 51.145 54.175 51.470 54.420 ;
        RECT 51.240 52.420 51.470 54.175 ;
        RECT 53.005 54.375 53.195 55.470 ;
        RECT 53.960 55.380 54.230 55.470 ;
        RECT 54.000 54.475 54.190 54.505 ;
        RECT 53.960 54.375 54.230 54.475 ;
        RECT 64.030 54.420 64.595 55.510 ;
        RECT 70.055 54.420 70.245 55.510 ;
        RECT 71.925 54.420 72.115 55.510 ;
        RECT 73.805 54.420 73.995 55.510 ;
        RECT 75.665 55.470 76.890 55.660 ;
        RECT 86.570 55.510 87.390 55.760 ;
        RECT 92.800 55.755 93.030 56.910 ;
        RECT 94.680 55.765 94.910 56.910 ;
        RECT 96.560 55.765 96.790 56.910 ;
        RECT 92.715 55.510 93.030 55.755 ;
        RECT 94.585 55.510 94.910 55.765 ;
        RECT 96.465 55.510 96.790 55.765 ;
        RECT 98.325 56.760 99.550 56.950 ;
        RECT 98.325 55.660 98.515 56.760 ;
        RECT 99.280 56.670 99.550 56.760 ;
        RECT 109.230 56.880 110.050 57.480 ;
        RECT 115.380 56.910 115.980 57.510 ;
        RECT 117.260 56.910 117.860 57.510 ;
        RECT 119.140 56.910 119.740 57.510 ;
        RECT 120.950 57.000 121.210 57.320 ;
        RECT 121.980 57.050 122.170 57.080 ;
        RECT 120.985 56.950 121.210 57.000 ;
        RECT 121.940 56.950 122.210 57.050 ;
        RECT 99.320 55.760 99.510 55.790 ;
        RECT 109.230 55.760 109.460 56.880 ;
        RECT 109.820 55.760 110.050 56.880 ;
        RECT 99.280 55.660 99.550 55.760 ;
        RECT 53.005 54.185 54.230 54.375 ;
        RECT 53.005 53.090 53.195 54.185 ;
        RECT 53.960 54.095 54.230 54.185 ;
        RECT 63.910 54.180 64.730 54.420 ;
        RECT 70.055 54.180 70.370 54.420 ;
        RECT 71.925 54.180 72.250 54.420 ;
        RECT 54.000 53.190 54.190 53.225 ;
        RECT 53.960 53.090 54.230 53.190 ;
        RECT 53.005 52.900 54.230 53.090 ;
        RECT 53.960 52.810 54.230 52.900 ;
        RECT 63.910 52.660 64.140 54.180 ;
        RECT 64.500 52.660 64.730 54.180 ;
        RECT 63.910 52.470 64.730 52.660 ;
        RECT 63.910 52.420 64.140 52.470 ;
        RECT 64.500 52.420 64.730 52.470 ;
        RECT 70.140 52.420 70.370 54.180 ;
        RECT 72.020 52.420 72.250 54.180 ;
        RECT 73.805 54.175 74.130 54.420 ;
        RECT 73.900 52.420 74.130 54.175 ;
        RECT 75.665 54.375 75.855 55.470 ;
        RECT 76.620 55.380 76.890 55.470 ;
        RECT 76.660 54.475 76.850 54.505 ;
        RECT 76.620 54.375 76.890 54.475 ;
        RECT 86.690 54.420 87.255 55.510 ;
        RECT 92.715 54.420 92.905 55.510 ;
        RECT 94.585 54.420 94.775 55.510 ;
        RECT 96.465 54.420 96.655 55.510 ;
        RECT 98.325 55.470 99.550 55.660 ;
        RECT 109.230 55.510 110.050 55.760 ;
        RECT 115.460 55.755 115.690 56.910 ;
        RECT 117.340 55.765 117.570 56.910 ;
        RECT 119.220 55.765 119.450 56.910 ;
        RECT 115.375 55.510 115.690 55.755 ;
        RECT 117.245 55.510 117.570 55.765 ;
        RECT 119.125 55.510 119.450 55.765 ;
        RECT 120.985 56.760 122.210 56.950 ;
        RECT 120.985 55.660 121.175 56.760 ;
        RECT 121.940 56.670 122.210 56.760 ;
        RECT 121.980 55.760 122.170 55.790 ;
        RECT 121.940 55.660 122.210 55.760 ;
        RECT 75.665 54.185 76.890 54.375 ;
        RECT 75.665 53.090 75.855 54.185 ;
        RECT 76.620 54.095 76.890 54.185 ;
        RECT 86.570 54.180 87.390 54.420 ;
        RECT 92.715 54.180 93.030 54.420 ;
        RECT 94.585 54.180 94.910 54.420 ;
        RECT 76.660 53.190 76.850 53.225 ;
        RECT 76.620 53.090 76.890 53.190 ;
        RECT 75.665 52.900 76.890 53.090 ;
        RECT 76.620 52.810 76.890 52.900 ;
        RECT 86.570 52.660 86.800 54.180 ;
        RECT 87.160 52.660 87.390 54.180 ;
        RECT 86.570 52.470 87.390 52.660 ;
        RECT 86.570 52.420 86.800 52.470 ;
        RECT 87.160 52.420 87.390 52.470 ;
        RECT 92.800 52.420 93.030 54.180 ;
        RECT 94.680 52.420 94.910 54.180 ;
        RECT 96.465 54.175 96.790 54.420 ;
        RECT 96.560 52.420 96.790 54.175 ;
        RECT 98.325 54.375 98.515 55.470 ;
        RECT 99.280 55.380 99.550 55.470 ;
        RECT 99.320 54.475 99.510 54.505 ;
        RECT 99.280 54.375 99.550 54.475 ;
        RECT 109.350 54.420 109.915 55.510 ;
        RECT 115.375 54.420 115.565 55.510 ;
        RECT 117.245 54.420 117.435 55.510 ;
        RECT 119.125 54.420 119.315 55.510 ;
        RECT 120.985 55.470 122.210 55.660 ;
        RECT 98.325 54.185 99.550 54.375 ;
        RECT 98.325 53.090 98.515 54.185 ;
        RECT 99.280 54.095 99.550 54.185 ;
        RECT 109.230 54.180 110.050 54.420 ;
        RECT 115.375 54.180 115.690 54.420 ;
        RECT 117.245 54.180 117.570 54.420 ;
        RECT 99.320 53.190 99.510 53.225 ;
        RECT 99.280 53.090 99.550 53.190 ;
        RECT 98.325 52.900 99.550 53.090 ;
        RECT 99.280 52.810 99.550 52.900 ;
        RECT 109.230 52.660 109.460 54.180 ;
        RECT 109.820 52.660 110.050 54.180 ;
        RECT 109.230 52.470 110.050 52.660 ;
        RECT 109.230 52.420 109.460 52.470 ;
        RECT 109.820 52.420 110.050 52.470 ;
        RECT 115.460 52.420 115.690 54.180 ;
        RECT 117.340 52.420 117.570 54.180 ;
        RECT 119.125 54.175 119.450 54.420 ;
        RECT 119.220 52.420 119.450 54.175 ;
        RECT 120.985 54.375 121.175 55.470 ;
        RECT 121.940 55.380 122.210 55.470 ;
        RECT 121.980 54.475 122.170 54.505 ;
        RECT 121.940 54.375 122.210 54.475 ;
        RECT 120.985 54.185 122.210 54.375 ;
        RECT 120.985 53.090 121.175 54.185 ;
        RECT 121.940 54.095 122.210 54.185 ;
        RECT 121.980 53.190 122.170 53.225 ;
        RECT 121.940 53.090 122.210 53.190 ;
        RECT 120.985 52.900 122.210 53.090 ;
        RECT 121.940 52.810 122.210 52.900 ;
      LAYER via ;
        RECT 59.520 183.740 59.780 184.000 ;
        RECT 59.840 183.740 60.100 184.000 ;
        RECT 60.160 183.740 60.420 184.000 ;
        RECT 60.480 183.740 60.740 184.000 ;
        RECT 60.800 183.740 61.060 184.000 ;
        RECT 78.030 183.740 78.290 184.000 ;
        RECT 78.350 183.740 78.610 184.000 ;
        RECT 78.670 183.740 78.930 184.000 ;
        RECT 78.990 183.740 79.250 184.000 ;
        RECT 79.310 183.740 79.570 184.000 ;
        RECT 96.540 183.740 96.800 184.000 ;
        RECT 96.860 183.740 97.120 184.000 ;
        RECT 97.180 183.740 97.440 184.000 ;
        RECT 97.500 183.740 97.760 184.000 ;
        RECT 97.820 183.740 98.080 184.000 ;
        RECT 115.050 183.740 115.310 184.000 ;
        RECT 115.370 183.740 115.630 184.000 ;
        RECT 115.690 183.740 115.950 184.000 ;
        RECT 116.010 183.740 116.270 184.000 ;
        RECT 116.330 183.740 116.590 184.000 ;
        RECT 59.520 178.300 59.780 178.560 ;
        RECT 59.840 178.300 60.100 178.560 ;
        RECT 60.160 178.300 60.420 178.560 ;
        RECT 60.480 178.300 60.740 178.560 ;
        RECT 60.800 178.300 61.060 178.560 ;
        RECT 78.030 178.300 78.290 178.560 ;
        RECT 78.350 178.300 78.610 178.560 ;
        RECT 78.670 178.300 78.930 178.560 ;
        RECT 78.990 178.300 79.250 178.560 ;
        RECT 79.310 178.300 79.570 178.560 ;
        RECT 96.540 178.300 96.800 178.560 ;
        RECT 96.860 178.300 97.120 178.560 ;
        RECT 97.180 178.300 97.440 178.560 ;
        RECT 97.500 178.300 97.760 178.560 ;
        RECT 97.820 178.300 98.080 178.560 ;
        RECT 115.050 178.300 115.310 178.560 ;
        RECT 115.370 178.300 115.630 178.560 ;
        RECT 115.690 178.300 115.950 178.560 ;
        RECT 116.010 178.300 116.270 178.560 ;
        RECT 116.330 178.300 116.590 178.560 ;
        RECT 59.520 172.860 59.780 173.120 ;
        RECT 59.840 172.860 60.100 173.120 ;
        RECT 60.160 172.860 60.420 173.120 ;
        RECT 60.480 172.860 60.740 173.120 ;
        RECT 60.800 172.860 61.060 173.120 ;
        RECT 78.030 172.860 78.290 173.120 ;
        RECT 78.350 172.860 78.610 173.120 ;
        RECT 78.670 172.860 78.930 173.120 ;
        RECT 78.990 172.860 79.250 173.120 ;
        RECT 79.310 172.860 79.570 173.120 ;
        RECT 96.540 172.860 96.800 173.120 ;
        RECT 96.860 172.860 97.120 173.120 ;
        RECT 97.180 172.860 97.440 173.120 ;
        RECT 97.500 172.860 97.760 173.120 ;
        RECT 97.820 172.860 98.080 173.120 ;
        RECT 115.050 172.860 115.310 173.120 ;
        RECT 115.370 172.860 115.630 173.120 ;
        RECT 115.690 172.860 115.950 173.120 ;
        RECT 116.010 172.860 116.270 173.120 ;
        RECT 116.330 172.860 116.590 173.120 ;
        RECT 59.520 167.420 59.780 167.680 ;
        RECT 59.840 167.420 60.100 167.680 ;
        RECT 60.160 167.420 60.420 167.680 ;
        RECT 60.480 167.420 60.740 167.680 ;
        RECT 60.800 167.420 61.060 167.680 ;
        RECT 78.030 167.420 78.290 167.680 ;
        RECT 78.350 167.420 78.610 167.680 ;
        RECT 78.670 167.420 78.930 167.680 ;
        RECT 78.990 167.420 79.250 167.680 ;
        RECT 79.310 167.420 79.570 167.680 ;
        RECT 96.540 167.420 96.800 167.680 ;
        RECT 96.860 167.420 97.120 167.680 ;
        RECT 97.180 167.420 97.440 167.680 ;
        RECT 97.500 167.420 97.760 167.680 ;
        RECT 97.820 167.420 98.080 167.680 ;
        RECT 115.050 167.420 115.310 167.680 ;
        RECT 115.370 167.420 115.630 167.680 ;
        RECT 115.690 167.420 115.950 167.680 ;
        RECT 116.010 167.420 116.270 167.680 ;
        RECT 116.330 167.420 116.590 167.680 ;
        RECT 59.520 161.980 59.780 162.240 ;
        RECT 59.840 161.980 60.100 162.240 ;
        RECT 60.160 161.980 60.420 162.240 ;
        RECT 60.480 161.980 60.740 162.240 ;
        RECT 60.800 161.980 61.060 162.240 ;
        RECT 78.030 161.980 78.290 162.240 ;
        RECT 78.350 161.980 78.610 162.240 ;
        RECT 78.670 161.980 78.930 162.240 ;
        RECT 78.990 161.980 79.250 162.240 ;
        RECT 79.310 161.980 79.570 162.240 ;
        RECT 96.540 161.980 96.800 162.240 ;
        RECT 96.860 161.980 97.120 162.240 ;
        RECT 97.180 161.980 97.440 162.240 ;
        RECT 97.500 161.980 97.760 162.240 ;
        RECT 97.820 161.980 98.080 162.240 ;
        RECT 115.050 161.980 115.310 162.240 ;
        RECT 115.370 161.980 115.630 162.240 ;
        RECT 115.690 161.980 115.950 162.240 ;
        RECT 116.010 161.980 116.270 162.240 ;
        RECT 116.330 161.980 116.590 162.240 ;
        RECT 59.520 156.540 59.780 156.800 ;
        RECT 59.840 156.540 60.100 156.800 ;
        RECT 60.160 156.540 60.420 156.800 ;
        RECT 60.480 156.540 60.740 156.800 ;
        RECT 60.800 156.540 61.060 156.800 ;
        RECT 78.030 156.540 78.290 156.800 ;
        RECT 78.350 156.540 78.610 156.800 ;
        RECT 78.670 156.540 78.930 156.800 ;
        RECT 78.990 156.540 79.250 156.800 ;
        RECT 79.310 156.540 79.570 156.800 ;
        RECT 96.540 156.540 96.800 156.800 ;
        RECT 96.860 156.540 97.120 156.800 ;
        RECT 97.180 156.540 97.440 156.800 ;
        RECT 97.500 156.540 97.760 156.800 ;
        RECT 97.820 156.540 98.080 156.800 ;
        RECT 115.050 156.540 115.310 156.800 ;
        RECT 115.370 156.540 115.630 156.800 ;
        RECT 115.690 156.540 115.950 156.800 ;
        RECT 116.010 156.540 116.270 156.800 ;
        RECT 116.330 156.540 116.590 156.800 ;
        RECT 63.940 126.930 64.700 127.470 ;
        RECT 70.090 126.960 70.630 127.500 ;
        RECT 71.970 126.960 72.510 127.500 ;
        RECT 73.850 126.960 74.390 127.500 ;
        RECT 75.630 127.050 75.890 127.310 ;
        RECT 86.600 126.930 87.360 127.470 ;
        RECT 92.750 126.960 93.290 127.500 ;
        RECT 94.630 126.960 95.170 127.500 ;
        RECT 96.510 126.960 97.050 127.500 ;
        RECT 98.290 127.050 98.550 127.310 ;
        RECT 109.260 126.930 110.020 127.470 ;
        RECT 115.410 126.960 115.950 127.500 ;
        RECT 117.290 126.960 117.830 127.500 ;
        RECT 119.170 126.960 119.710 127.500 ;
        RECT 120.950 127.050 121.210 127.310 ;
        RECT 61.290 121.620 62.210 122.540 ;
        RECT 83.950 121.620 84.870 122.540 ;
        RECT 106.610 121.620 107.530 122.540 ;
        RECT 124.200 124.620 124.550 126.780 ;
        RECT 41.280 109.590 42.040 110.130 ;
        RECT 47.430 109.620 47.970 110.160 ;
        RECT 49.310 109.620 49.850 110.160 ;
        RECT 51.190 109.620 51.730 110.160 ;
        RECT 52.970 109.710 53.230 109.970 ;
        RECT 63.940 109.590 64.700 110.130 ;
        RECT 70.090 109.620 70.630 110.160 ;
        RECT 71.970 109.620 72.510 110.160 ;
        RECT 73.850 109.620 74.390 110.160 ;
        RECT 75.630 109.710 75.890 109.970 ;
        RECT 86.600 109.590 87.360 110.130 ;
        RECT 92.750 109.620 93.290 110.160 ;
        RECT 94.630 109.620 95.170 110.160 ;
        RECT 96.510 109.620 97.050 110.160 ;
        RECT 98.290 109.710 98.550 109.970 ;
        RECT 38.630 104.280 39.550 105.200 ;
        RECT 109.260 109.590 110.020 110.130 ;
        RECT 115.410 109.620 115.950 110.160 ;
        RECT 117.290 109.620 117.830 110.160 ;
        RECT 119.170 109.620 119.710 110.160 ;
        RECT 120.950 109.710 121.210 109.970 ;
        RECT 61.290 104.280 62.210 105.200 ;
        RECT 83.950 104.280 84.870 105.200 ;
        RECT 106.610 104.280 107.530 105.200 ;
        RECT 41.280 92.250 42.040 92.790 ;
        RECT 47.430 92.280 47.970 92.820 ;
        RECT 49.310 92.280 49.850 92.820 ;
        RECT 51.190 92.280 51.730 92.820 ;
        RECT 52.970 92.370 53.230 92.630 ;
        RECT 63.940 92.250 64.700 92.790 ;
        RECT 70.090 92.280 70.630 92.820 ;
        RECT 71.970 92.280 72.510 92.820 ;
        RECT 73.850 92.280 74.390 92.820 ;
        RECT 75.630 92.370 75.890 92.630 ;
        RECT 86.600 92.250 87.360 92.790 ;
        RECT 92.750 92.280 93.290 92.820 ;
        RECT 94.630 92.280 95.170 92.820 ;
        RECT 96.510 92.280 97.050 92.820 ;
        RECT 98.290 92.370 98.550 92.630 ;
        RECT 38.630 86.940 39.550 87.860 ;
        RECT 109.260 92.250 110.020 92.790 ;
        RECT 115.410 92.280 115.950 92.820 ;
        RECT 117.290 92.280 117.830 92.820 ;
        RECT 119.170 92.280 119.710 92.820 ;
        RECT 120.950 92.370 121.210 92.630 ;
        RECT 61.290 86.940 62.210 87.860 ;
        RECT 83.950 86.940 84.870 87.860 ;
        RECT 106.610 86.940 107.530 87.860 ;
        RECT 41.280 74.910 42.040 75.450 ;
        RECT 47.430 74.940 47.970 75.480 ;
        RECT 49.310 74.940 49.850 75.480 ;
        RECT 51.190 74.940 51.730 75.480 ;
        RECT 52.970 75.030 53.230 75.290 ;
        RECT 63.940 74.910 64.700 75.450 ;
        RECT 70.090 74.940 70.630 75.480 ;
        RECT 71.970 74.940 72.510 75.480 ;
        RECT 73.850 74.940 74.390 75.480 ;
        RECT 75.630 75.030 75.890 75.290 ;
        RECT 86.600 74.910 87.360 75.450 ;
        RECT 92.750 74.940 93.290 75.480 ;
        RECT 94.630 74.940 95.170 75.480 ;
        RECT 96.510 74.940 97.050 75.480 ;
        RECT 98.290 75.030 98.550 75.290 ;
        RECT 38.630 69.600 39.550 70.520 ;
        RECT 109.260 74.910 110.020 75.450 ;
        RECT 115.410 74.940 115.950 75.480 ;
        RECT 117.290 74.940 117.830 75.480 ;
        RECT 119.170 74.940 119.710 75.480 ;
        RECT 120.950 75.030 121.210 75.290 ;
        RECT 61.290 69.600 62.210 70.520 ;
        RECT 83.950 69.600 84.870 70.520 ;
        RECT 106.610 69.600 107.530 70.520 ;
        RECT 41.280 56.910 42.040 57.450 ;
        RECT 47.430 56.940 47.970 57.480 ;
        RECT 49.310 56.940 49.850 57.480 ;
        RECT 51.190 56.940 51.730 57.480 ;
        RECT 52.970 57.030 53.230 57.290 ;
        RECT 63.940 56.910 64.700 57.450 ;
        RECT 70.090 56.940 70.630 57.480 ;
        RECT 71.970 56.940 72.510 57.480 ;
        RECT 73.850 56.940 74.390 57.480 ;
        RECT 75.630 57.030 75.890 57.290 ;
        RECT 86.600 56.910 87.360 57.450 ;
        RECT 92.750 56.940 93.290 57.480 ;
        RECT 94.630 56.940 95.170 57.480 ;
        RECT 96.510 56.940 97.050 57.480 ;
        RECT 98.290 57.030 98.550 57.290 ;
        RECT 109.260 56.910 110.020 57.450 ;
        RECT 115.410 56.940 115.950 57.480 ;
        RECT 117.290 56.940 117.830 57.480 ;
        RECT 119.170 56.940 119.710 57.480 ;
        RECT 120.950 57.030 121.210 57.290 ;
      LAYER met2 ;
        RECT 59.520 183.685 61.060 184.055 ;
        RECT 78.030 183.685 79.570 184.055 ;
        RECT 96.540 183.685 98.080 184.055 ;
        RECT 115.050 183.685 116.590 184.055 ;
        RECT 59.520 178.245 61.060 178.615 ;
        RECT 78.030 178.245 79.570 178.615 ;
        RECT 96.540 178.245 98.080 178.615 ;
        RECT 115.050 178.245 116.590 178.615 ;
        RECT 59.520 172.805 61.060 173.175 ;
        RECT 78.030 172.805 79.570 173.175 ;
        RECT 96.540 172.805 98.080 173.175 ;
        RECT 115.050 172.805 116.590 173.175 ;
        RECT 59.520 167.365 61.060 167.735 ;
        RECT 78.030 167.365 79.570 167.735 ;
        RECT 96.540 167.365 98.080 167.735 ;
        RECT 115.050 167.365 116.590 167.735 ;
        RECT 59.520 161.925 61.060 162.295 ;
        RECT 78.030 161.925 79.570 162.295 ;
        RECT 96.540 161.925 98.080 162.295 ;
        RECT 115.050 161.925 116.590 162.295 ;
        RECT 59.520 156.485 61.060 156.855 ;
        RECT 78.030 156.485 79.570 156.855 ;
        RECT 96.540 156.485 98.080 156.855 ;
        RECT 115.050 156.485 116.590 156.855 ;
        RECT 63.670 127.320 64.990 127.510 ;
        RECT 69.710 127.320 71.030 127.530 ;
        RECT 71.590 127.320 72.910 127.530 ;
        RECT 73.470 127.320 74.790 127.540 ;
        RECT 75.890 127.320 76.890 128.010 ;
        RECT 86.330 127.320 87.650 127.510 ;
        RECT 92.370 127.320 93.690 127.530 ;
        RECT 94.250 127.320 95.570 127.530 ;
        RECT 96.130 127.320 97.450 127.540 ;
        RECT 98.550 127.320 99.550 128.010 ;
        RECT 108.990 127.320 110.310 127.510 ;
        RECT 115.030 127.320 116.350 127.530 ;
        RECT 116.910 127.320 118.230 127.530 ;
        RECT 118.790 127.320 120.110 127.540 ;
        RECT 121.210 127.320 122.210 128.010 ;
        RECT 123.875 127.810 124.875 128.810 ;
        RECT 62.480 127.080 76.890 127.320 ;
        RECT 30.920 55.395 31.920 125.475 ;
        RECT 62.480 123.470 62.720 127.080 ;
        RECT 63.670 126.750 64.990 127.080 ;
        RECT 69.710 126.770 71.030 127.080 ;
        RECT 71.590 126.770 72.910 127.080 ;
        RECT 73.470 126.780 74.790 127.080 ;
        RECT 75.600 127.050 76.890 127.080 ;
        RECT 75.890 127.010 76.890 127.050 ;
        RECT 85.140 127.080 99.550 127.320 ;
        RECT 85.140 123.470 85.380 127.080 ;
        RECT 86.330 126.750 87.650 127.080 ;
        RECT 92.370 126.770 93.690 127.080 ;
        RECT 94.250 126.770 95.570 127.080 ;
        RECT 96.130 126.780 97.450 127.080 ;
        RECT 98.260 127.050 99.550 127.080 ;
        RECT 98.550 127.010 99.550 127.050 ;
        RECT 107.800 127.080 122.210 127.320 ;
        RECT 107.800 123.470 108.040 127.080 ;
        RECT 108.990 126.750 110.310 127.080 ;
        RECT 115.030 126.770 116.350 127.080 ;
        RECT 116.910 126.770 118.230 127.080 ;
        RECT 118.790 126.780 120.110 127.080 ;
        RECT 120.920 127.050 122.210 127.080 ;
        RECT 121.210 127.010 122.210 127.050 ;
        RECT 124.250 126.810 124.500 127.810 ;
        RECT 124.200 124.590 124.550 126.810 ;
        RECT 61.960 123.230 62.720 123.470 ;
        RECT 84.620 123.230 85.380 123.470 ;
        RECT 107.280 123.230 108.040 123.470 ;
        RECT 61.960 122.580 62.200 123.230 ;
        RECT 84.620 122.580 84.860 123.230 ;
        RECT 107.280 122.580 107.520 123.230 ;
        RECT 61.250 121.580 62.250 122.580 ;
        RECT 83.910 121.580 84.910 122.580 ;
        RECT 106.570 121.580 107.570 122.580 ;
        RECT 41.010 109.980 42.330 110.170 ;
        RECT 47.050 109.980 48.370 110.190 ;
        RECT 48.930 109.980 50.250 110.190 ;
        RECT 50.810 109.980 52.130 110.200 ;
        RECT 53.230 109.980 54.230 110.670 ;
        RECT 63.670 109.980 64.990 110.170 ;
        RECT 69.710 109.980 71.030 110.190 ;
        RECT 71.590 109.980 72.910 110.190 ;
        RECT 73.470 109.980 74.790 110.200 ;
        RECT 75.890 109.980 76.890 110.670 ;
        RECT 86.330 109.980 87.650 110.170 ;
        RECT 92.370 109.980 93.690 110.190 ;
        RECT 94.250 109.980 95.570 110.190 ;
        RECT 96.130 109.980 97.450 110.200 ;
        RECT 98.550 109.980 99.550 110.670 ;
        RECT 108.990 109.980 110.310 110.170 ;
        RECT 115.030 109.980 116.350 110.190 ;
        RECT 116.910 109.980 118.230 110.190 ;
        RECT 118.790 109.980 120.110 110.200 ;
        RECT 121.210 109.980 122.210 110.670 ;
        RECT 39.820 109.740 54.230 109.980 ;
        RECT 39.820 106.130 40.060 109.740 ;
        RECT 41.010 109.410 42.330 109.740 ;
        RECT 47.050 109.430 48.370 109.740 ;
        RECT 48.930 109.430 50.250 109.740 ;
        RECT 50.810 109.440 52.130 109.740 ;
        RECT 52.940 109.710 54.230 109.740 ;
        RECT 53.230 109.670 54.230 109.710 ;
        RECT 62.480 109.740 76.890 109.980 ;
        RECT 62.480 106.130 62.720 109.740 ;
        RECT 63.670 109.410 64.990 109.740 ;
        RECT 69.710 109.430 71.030 109.740 ;
        RECT 71.590 109.430 72.910 109.740 ;
        RECT 73.470 109.440 74.790 109.740 ;
        RECT 75.600 109.710 76.890 109.740 ;
        RECT 75.890 109.670 76.890 109.710 ;
        RECT 85.140 109.740 99.550 109.980 ;
        RECT 85.140 106.130 85.380 109.740 ;
        RECT 86.330 109.410 87.650 109.740 ;
        RECT 92.370 109.430 93.690 109.740 ;
        RECT 94.250 109.430 95.570 109.740 ;
        RECT 96.130 109.440 97.450 109.740 ;
        RECT 98.260 109.710 99.550 109.740 ;
        RECT 98.550 109.670 99.550 109.710 ;
        RECT 107.800 109.740 122.210 109.980 ;
        RECT 107.800 106.130 108.040 109.740 ;
        RECT 108.990 109.410 110.310 109.740 ;
        RECT 115.030 109.430 116.350 109.740 ;
        RECT 116.910 109.430 118.230 109.740 ;
        RECT 118.790 109.440 120.110 109.740 ;
        RECT 120.920 109.710 122.210 109.740 ;
        RECT 121.210 109.670 122.210 109.710 ;
        RECT 39.300 105.890 40.060 106.130 ;
        RECT 61.960 105.890 62.720 106.130 ;
        RECT 84.620 105.890 85.380 106.130 ;
        RECT 107.280 105.890 108.040 106.130 ;
        RECT 39.300 105.240 39.540 105.890 ;
        RECT 61.960 105.240 62.200 105.890 ;
        RECT 84.620 105.240 84.860 105.890 ;
        RECT 107.280 105.240 107.520 105.890 ;
        RECT 38.590 104.240 39.590 105.240 ;
        RECT 61.250 104.240 62.250 105.240 ;
        RECT 83.910 104.240 84.910 105.240 ;
        RECT 106.570 104.240 107.570 105.240 ;
        RECT 41.010 92.640 42.330 92.830 ;
        RECT 47.050 92.640 48.370 92.850 ;
        RECT 48.930 92.640 50.250 92.850 ;
        RECT 50.810 92.640 52.130 92.860 ;
        RECT 53.230 92.640 54.230 93.330 ;
        RECT 63.670 92.640 64.990 92.830 ;
        RECT 69.710 92.640 71.030 92.850 ;
        RECT 71.590 92.640 72.910 92.850 ;
        RECT 73.470 92.640 74.790 92.860 ;
        RECT 75.890 92.640 76.890 93.330 ;
        RECT 86.330 92.640 87.650 92.830 ;
        RECT 92.370 92.640 93.690 92.850 ;
        RECT 94.250 92.640 95.570 92.850 ;
        RECT 96.130 92.640 97.450 92.860 ;
        RECT 98.550 92.640 99.550 93.330 ;
        RECT 108.990 92.640 110.310 92.830 ;
        RECT 115.030 92.640 116.350 92.850 ;
        RECT 116.910 92.640 118.230 92.850 ;
        RECT 118.790 92.640 120.110 92.860 ;
        RECT 121.210 92.640 122.210 93.330 ;
        RECT 39.820 92.400 54.230 92.640 ;
        RECT 39.820 88.790 40.060 92.400 ;
        RECT 41.010 92.070 42.330 92.400 ;
        RECT 47.050 92.090 48.370 92.400 ;
        RECT 48.930 92.090 50.250 92.400 ;
        RECT 50.810 92.100 52.130 92.400 ;
        RECT 52.940 92.370 54.230 92.400 ;
        RECT 53.230 92.330 54.230 92.370 ;
        RECT 62.480 92.400 76.890 92.640 ;
        RECT 62.480 88.790 62.720 92.400 ;
        RECT 63.670 92.070 64.990 92.400 ;
        RECT 69.710 92.090 71.030 92.400 ;
        RECT 71.590 92.090 72.910 92.400 ;
        RECT 73.470 92.100 74.790 92.400 ;
        RECT 75.600 92.370 76.890 92.400 ;
        RECT 75.890 92.330 76.890 92.370 ;
        RECT 85.140 92.400 99.550 92.640 ;
        RECT 85.140 88.790 85.380 92.400 ;
        RECT 86.330 92.070 87.650 92.400 ;
        RECT 92.370 92.090 93.690 92.400 ;
        RECT 94.250 92.090 95.570 92.400 ;
        RECT 96.130 92.100 97.450 92.400 ;
        RECT 98.260 92.370 99.550 92.400 ;
        RECT 98.550 92.330 99.550 92.370 ;
        RECT 107.800 92.400 122.210 92.640 ;
        RECT 107.800 88.790 108.040 92.400 ;
        RECT 108.990 92.070 110.310 92.400 ;
        RECT 115.030 92.090 116.350 92.400 ;
        RECT 116.910 92.090 118.230 92.400 ;
        RECT 118.790 92.100 120.110 92.400 ;
        RECT 120.920 92.370 122.210 92.400 ;
        RECT 121.210 92.330 122.210 92.370 ;
        RECT 39.300 88.550 40.060 88.790 ;
        RECT 61.960 88.550 62.720 88.790 ;
        RECT 84.620 88.550 85.380 88.790 ;
        RECT 107.280 88.550 108.040 88.790 ;
        RECT 39.300 87.900 39.540 88.550 ;
        RECT 61.960 87.900 62.200 88.550 ;
        RECT 84.620 87.900 84.860 88.550 ;
        RECT 107.280 87.900 107.520 88.550 ;
        RECT 38.590 86.900 39.590 87.900 ;
        RECT 61.250 86.900 62.250 87.900 ;
        RECT 83.910 86.900 84.910 87.900 ;
        RECT 106.570 86.900 107.570 87.900 ;
        RECT 41.010 75.300 42.330 75.490 ;
        RECT 47.050 75.300 48.370 75.510 ;
        RECT 48.930 75.300 50.250 75.510 ;
        RECT 50.810 75.300 52.130 75.520 ;
        RECT 53.230 75.300 54.230 75.990 ;
        RECT 63.670 75.300 64.990 75.490 ;
        RECT 69.710 75.300 71.030 75.510 ;
        RECT 71.590 75.300 72.910 75.510 ;
        RECT 73.470 75.300 74.790 75.520 ;
        RECT 75.890 75.300 76.890 75.990 ;
        RECT 86.330 75.300 87.650 75.490 ;
        RECT 92.370 75.300 93.690 75.510 ;
        RECT 94.250 75.300 95.570 75.510 ;
        RECT 96.130 75.300 97.450 75.520 ;
        RECT 98.550 75.300 99.550 75.990 ;
        RECT 108.990 75.300 110.310 75.490 ;
        RECT 115.030 75.300 116.350 75.510 ;
        RECT 116.910 75.300 118.230 75.510 ;
        RECT 118.790 75.300 120.110 75.520 ;
        RECT 121.210 75.300 122.210 75.990 ;
        RECT 39.820 75.060 54.230 75.300 ;
        RECT 39.820 71.450 40.060 75.060 ;
        RECT 41.010 74.730 42.330 75.060 ;
        RECT 47.050 74.750 48.370 75.060 ;
        RECT 48.930 74.750 50.250 75.060 ;
        RECT 50.810 74.760 52.130 75.060 ;
        RECT 52.940 75.030 54.230 75.060 ;
        RECT 53.230 74.990 54.230 75.030 ;
        RECT 62.480 75.060 76.890 75.300 ;
        RECT 62.480 71.450 62.720 75.060 ;
        RECT 63.670 74.730 64.990 75.060 ;
        RECT 69.710 74.750 71.030 75.060 ;
        RECT 71.590 74.750 72.910 75.060 ;
        RECT 73.470 74.760 74.790 75.060 ;
        RECT 75.600 75.030 76.890 75.060 ;
        RECT 75.890 74.990 76.890 75.030 ;
        RECT 85.140 75.060 99.550 75.300 ;
        RECT 85.140 71.450 85.380 75.060 ;
        RECT 86.330 74.730 87.650 75.060 ;
        RECT 92.370 74.750 93.690 75.060 ;
        RECT 94.250 74.750 95.570 75.060 ;
        RECT 96.130 74.760 97.450 75.060 ;
        RECT 98.260 75.030 99.550 75.060 ;
        RECT 98.550 74.990 99.550 75.030 ;
        RECT 107.800 75.060 122.210 75.300 ;
        RECT 107.800 71.450 108.040 75.060 ;
        RECT 108.990 74.730 110.310 75.060 ;
        RECT 115.030 74.750 116.350 75.060 ;
        RECT 116.910 74.750 118.230 75.060 ;
        RECT 118.790 74.760 120.110 75.060 ;
        RECT 120.920 75.030 122.210 75.060 ;
        RECT 121.210 74.990 122.210 75.030 ;
        RECT 39.300 71.210 40.060 71.450 ;
        RECT 61.960 71.210 62.720 71.450 ;
        RECT 84.620 71.210 85.380 71.450 ;
        RECT 107.280 71.210 108.040 71.450 ;
        RECT 39.300 70.560 39.540 71.210 ;
        RECT 61.960 70.560 62.200 71.210 ;
        RECT 84.620 70.560 84.860 71.210 ;
        RECT 107.280 70.560 107.520 71.210 ;
        RECT 38.590 69.560 39.590 70.560 ;
        RECT 61.250 69.560 62.250 70.560 ;
        RECT 83.910 69.560 84.910 70.560 ;
        RECT 106.570 69.560 107.570 70.560 ;
        RECT 41.010 57.300 42.330 57.490 ;
        RECT 47.050 57.300 48.370 57.510 ;
        RECT 48.930 57.300 50.250 57.510 ;
        RECT 50.810 57.300 52.130 57.520 ;
        RECT 53.230 57.300 54.230 57.990 ;
        RECT 41.010 57.060 54.230 57.300 ;
        RECT 41.010 56.730 42.330 57.060 ;
        RECT 47.050 56.750 48.370 57.060 ;
        RECT 48.930 56.750 50.250 57.060 ;
        RECT 50.810 56.760 52.130 57.060 ;
        RECT 52.940 57.030 54.230 57.060 ;
        RECT 53.230 56.990 54.230 57.030 ;
        RECT 63.670 57.300 64.990 57.490 ;
        RECT 69.710 57.300 71.030 57.510 ;
        RECT 71.590 57.300 72.910 57.510 ;
        RECT 73.470 57.300 74.790 57.520 ;
        RECT 75.890 57.300 76.890 57.990 ;
        RECT 63.670 57.060 76.890 57.300 ;
        RECT 63.670 56.730 64.990 57.060 ;
        RECT 69.710 56.750 71.030 57.060 ;
        RECT 71.590 56.750 72.910 57.060 ;
        RECT 73.470 56.760 74.790 57.060 ;
        RECT 75.600 57.030 76.890 57.060 ;
        RECT 75.890 56.990 76.890 57.030 ;
        RECT 86.330 57.300 87.650 57.490 ;
        RECT 92.370 57.300 93.690 57.510 ;
        RECT 94.250 57.300 95.570 57.510 ;
        RECT 96.130 57.300 97.450 57.520 ;
        RECT 98.550 57.300 99.550 57.990 ;
        RECT 86.330 57.060 99.550 57.300 ;
        RECT 86.330 56.730 87.650 57.060 ;
        RECT 92.370 56.750 93.690 57.060 ;
        RECT 94.250 56.750 95.570 57.060 ;
        RECT 96.130 56.760 97.450 57.060 ;
        RECT 98.260 57.030 99.550 57.060 ;
        RECT 98.550 56.990 99.550 57.030 ;
        RECT 108.990 57.300 110.310 57.490 ;
        RECT 115.030 57.300 116.350 57.510 ;
        RECT 116.910 57.300 118.230 57.510 ;
        RECT 118.790 57.300 120.110 57.520 ;
        RECT 121.210 57.300 122.210 57.990 ;
        RECT 108.990 57.060 122.210 57.300 ;
        RECT 108.990 56.730 110.310 57.060 ;
        RECT 115.030 56.750 116.350 57.060 ;
        RECT 116.910 56.750 118.230 57.060 ;
        RECT 118.790 56.760 120.110 57.060 ;
        RECT 120.920 57.030 122.210 57.060 ;
        RECT 121.210 56.990 122.210 57.030 ;
        RECT 30.900 54.445 31.940 55.395 ;
        RECT 30.920 54.420 31.920 54.445 ;
        RECT 127.800 54.385 128.800 125.485 ;
      LAYER via2 ;
        RECT 59.550 183.730 59.830 184.010 ;
        RECT 59.950 183.730 60.230 184.010 ;
        RECT 60.350 183.730 60.630 184.010 ;
        RECT 60.750 183.730 61.030 184.010 ;
        RECT 78.060 183.730 78.340 184.010 ;
        RECT 78.460 183.730 78.740 184.010 ;
        RECT 78.860 183.730 79.140 184.010 ;
        RECT 79.260 183.730 79.540 184.010 ;
        RECT 96.570 183.730 96.850 184.010 ;
        RECT 96.970 183.730 97.250 184.010 ;
        RECT 97.370 183.730 97.650 184.010 ;
        RECT 97.770 183.730 98.050 184.010 ;
        RECT 115.080 183.730 115.360 184.010 ;
        RECT 115.480 183.730 115.760 184.010 ;
        RECT 115.880 183.730 116.160 184.010 ;
        RECT 116.280 183.730 116.560 184.010 ;
        RECT 59.550 178.290 59.830 178.570 ;
        RECT 59.950 178.290 60.230 178.570 ;
        RECT 60.350 178.290 60.630 178.570 ;
        RECT 60.750 178.290 61.030 178.570 ;
        RECT 78.060 178.290 78.340 178.570 ;
        RECT 78.460 178.290 78.740 178.570 ;
        RECT 78.860 178.290 79.140 178.570 ;
        RECT 79.260 178.290 79.540 178.570 ;
        RECT 96.570 178.290 96.850 178.570 ;
        RECT 96.970 178.290 97.250 178.570 ;
        RECT 97.370 178.290 97.650 178.570 ;
        RECT 97.770 178.290 98.050 178.570 ;
        RECT 115.080 178.290 115.360 178.570 ;
        RECT 115.480 178.290 115.760 178.570 ;
        RECT 115.880 178.290 116.160 178.570 ;
        RECT 116.280 178.290 116.560 178.570 ;
        RECT 59.550 172.850 59.830 173.130 ;
        RECT 59.950 172.850 60.230 173.130 ;
        RECT 60.350 172.850 60.630 173.130 ;
        RECT 60.750 172.850 61.030 173.130 ;
        RECT 78.060 172.850 78.340 173.130 ;
        RECT 78.460 172.850 78.740 173.130 ;
        RECT 78.860 172.850 79.140 173.130 ;
        RECT 79.260 172.850 79.540 173.130 ;
        RECT 96.570 172.850 96.850 173.130 ;
        RECT 96.970 172.850 97.250 173.130 ;
        RECT 97.370 172.850 97.650 173.130 ;
        RECT 97.770 172.850 98.050 173.130 ;
        RECT 115.080 172.850 115.360 173.130 ;
        RECT 115.480 172.850 115.760 173.130 ;
        RECT 115.880 172.850 116.160 173.130 ;
        RECT 116.280 172.850 116.560 173.130 ;
        RECT 59.550 167.410 59.830 167.690 ;
        RECT 59.950 167.410 60.230 167.690 ;
        RECT 60.350 167.410 60.630 167.690 ;
        RECT 60.750 167.410 61.030 167.690 ;
        RECT 78.060 167.410 78.340 167.690 ;
        RECT 78.460 167.410 78.740 167.690 ;
        RECT 78.860 167.410 79.140 167.690 ;
        RECT 79.260 167.410 79.540 167.690 ;
        RECT 96.570 167.410 96.850 167.690 ;
        RECT 96.970 167.410 97.250 167.690 ;
        RECT 97.370 167.410 97.650 167.690 ;
        RECT 97.770 167.410 98.050 167.690 ;
        RECT 115.080 167.410 115.360 167.690 ;
        RECT 115.480 167.410 115.760 167.690 ;
        RECT 115.880 167.410 116.160 167.690 ;
        RECT 116.280 167.410 116.560 167.690 ;
        RECT 59.550 161.970 59.830 162.250 ;
        RECT 59.950 161.970 60.230 162.250 ;
        RECT 60.350 161.970 60.630 162.250 ;
        RECT 60.750 161.970 61.030 162.250 ;
        RECT 78.060 161.970 78.340 162.250 ;
        RECT 78.460 161.970 78.740 162.250 ;
        RECT 78.860 161.970 79.140 162.250 ;
        RECT 79.260 161.970 79.540 162.250 ;
        RECT 96.570 161.970 96.850 162.250 ;
        RECT 96.970 161.970 97.250 162.250 ;
        RECT 97.370 161.970 97.650 162.250 ;
        RECT 97.770 161.970 98.050 162.250 ;
        RECT 115.080 161.970 115.360 162.250 ;
        RECT 115.480 161.970 115.760 162.250 ;
        RECT 115.880 161.970 116.160 162.250 ;
        RECT 116.280 161.970 116.560 162.250 ;
        RECT 59.550 156.530 59.830 156.810 ;
        RECT 59.950 156.530 60.230 156.810 ;
        RECT 60.350 156.530 60.630 156.810 ;
        RECT 60.750 156.530 61.030 156.810 ;
        RECT 78.060 156.530 78.340 156.810 ;
        RECT 78.460 156.530 78.740 156.810 ;
        RECT 78.860 156.530 79.140 156.810 ;
        RECT 79.260 156.530 79.540 156.810 ;
        RECT 96.570 156.530 96.850 156.810 ;
        RECT 96.970 156.530 97.250 156.810 ;
        RECT 97.370 156.530 97.650 156.810 ;
        RECT 97.770 156.530 98.050 156.810 ;
        RECT 115.080 156.530 115.360 156.810 ;
        RECT 115.480 156.530 115.760 156.810 ;
        RECT 115.880 156.530 116.160 156.810 ;
        RECT 116.280 156.530 116.560 156.810 ;
        RECT 30.920 124.430 31.920 125.430 ;
        RECT 63.720 126.800 64.940 127.460 ;
        RECT 69.760 126.820 70.980 127.480 ;
        RECT 71.640 126.820 72.860 127.480 ;
        RECT 73.520 126.830 74.740 127.490 ;
        RECT 75.940 127.060 76.840 127.960 ;
        RECT 86.380 126.800 87.600 127.460 ;
        RECT 92.420 126.820 93.640 127.480 ;
        RECT 94.300 126.820 95.520 127.480 ;
        RECT 96.180 126.830 97.400 127.490 ;
        RECT 98.600 127.060 99.500 127.960 ;
        RECT 109.040 126.800 110.260 127.460 ;
        RECT 115.080 126.820 116.300 127.480 ;
        RECT 116.960 126.820 118.180 127.480 ;
        RECT 118.840 126.830 120.060 127.490 ;
        RECT 121.260 127.060 122.160 127.960 ;
        RECT 123.925 127.860 124.825 128.760 ;
        RECT 127.800 124.440 128.800 125.440 ;
        RECT 61.300 121.630 62.200 122.530 ;
        RECT 83.960 121.630 84.860 122.530 ;
        RECT 106.620 121.630 107.520 122.530 ;
        RECT 30.920 107.120 31.920 108.120 ;
        RECT 41.060 109.460 42.280 110.120 ;
        RECT 47.100 109.480 48.320 110.140 ;
        RECT 48.980 109.480 50.200 110.140 ;
        RECT 50.860 109.490 52.080 110.150 ;
        RECT 53.280 109.720 54.180 110.620 ;
        RECT 63.720 109.460 64.940 110.120 ;
        RECT 69.760 109.480 70.980 110.140 ;
        RECT 71.640 109.480 72.860 110.140 ;
        RECT 73.520 109.490 74.740 110.150 ;
        RECT 75.940 109.720 76.840 110.620 ;
        RECT 86.380 109.460 87.600 110.120 ;
        RECT 92.420 109.480 93.640 110.140 ;
        RECT 94.300 109.480 95.520 110.140 ;
        RECT 96.180 109.490 97.400 110.150 ;
        RECT 98.600 109.720 99.500 110.620 ;
        RECT 109.040 109.460 110.260 110.120 ;
        RECT 115.080 109.480 116.300 110.140 ;
        RECT 116.960 109.480 118.180 110.140 ;
        RECT 118.840 109.490 120.060 110.150 ;
        RECT 121.260 109.720 122.160 110.620 ;
        RECT 127.800 107.100 128.800 108.100 ;
        RECT 38.640 104.290 39.540 105.190 ;
        RECT 61.300 104.290 62.200 105.190 ;
        RECT 83.960 104.290 84.860 105.190 ;
        RECT 106.620 104.290 107.520 105.190 ;
        RECT 30.920 89.760 31.920 90.760 ;
        RECT 41.060 92.120 42.280 92.780 ;
        RECT 47.100 92.140 48.320 92.800 ;
        RECT 48.980 92.140 50.200 92.800 ;
        RECT 50.860 92.150 52.080 92.810 ;
        RECT 53.280 92.380 54.180 93.280 ;
        RECT 63.720 92.120 64.940 92.780 ;
        RECT 69.760 92.140 70.980 92.800 ;
        RECT 71.640 92.140 72.860 92.800 ;
        RECT 73.520 92.150 74.740 92.810 ;
        RECT 75.940 92.380 76.840 93.280 ;
        RECT 86.380 92.120 87.600 92.780 ;
        RECT 92.420 92.140 93.640 92.800 ;
        RECT 94.300 92.140 95.520 92.800 ;
        RECT 96.180 92.150 97.400 92.810 ;
        RECT 98.600 92.380 99.500 93.280 ;
        RECT 109.040 92.120 110.260 92.780 ;
        RECT 115.080 92.140 116.300 92.800 ;
        RECT 116.960 92.140 118.180 92.800 ;
        RECT 118.840 92.150 120.060 92.810 ;
        RECT 121.260 92.380 122.160 93.280 ;
        RECT 127.800 89.750 128.800 90.750 ;
        RECT 38.640 86.950 39.540 87.850 ;
        RECT 61.300 86.950 62.200 87.850 ;
        RECT 83.960 86.950 84.860 87.850 ;
        RECT 106.620 86.950 107.520 87.850 ;
        RECT 30.920 72.440 31.920 73.440 ;
        RECT 41.060 74.780 42.280 75.440 ;
        RECT 47.100 74.800 48.320 75.460 ;
        RECT 48.980 74.800 50.200 75.460 ;
        RECT 50.860 74.810 52.080 75.470 ;
        RECT 53.280 75.040 54.180 75.940 ;
        RECT 63.720 74.780 64.940 75.440 ;
        RECT 69.760 74.800 70.980 75.460 ;
        RECT 71.640 74.800 72.860 75.460 ;
        RECT 73.520 74.810 74.740 75.470 ;
        RECT 75.940 75.040 76.840 75.940 ;
        RECT 86.380 74.780 87.600 75.440 ;
        RECT 92.420 74.800 93.640 75.460 ;
        RECT 94.300 74.800 95.520 75.460 ;
        RECT 96.180 74.810 97.400 75.470 ;
        RECT 98.600 75.040 99.500 75.940 ;
        RECT 109.040 74.780 110.260 75.440 ;
        RECT 115.080 74.800 116.300 75.460 ;
        RECT 116.960 74.800 118.180 75.460 ;
        RECT 118.840 74.810 120.060 75.470 ;
        RECT 121.260 75.040 122.160 75.940 ;
        RECT 127.800 72.420 128.800 73.420 ;
        RECT 38.640 69.610 39.540 70.510 ;
        RECT 61.300 69.610 62.200 70.510 ;
        RECT 83.960 69.610 84.860 70.510 ;
        RECT 106.620 69.610 107.520 70.510 ;
        RECT 41.060 56.780 42.280 57.440 ;
        RECT 47.100 56.800 48.320 57.460 ;
        RECT 48.980 56.800 50.200 57.460 ;
        RECT 50.860 56.810 52.080 57.470 ;
        RECT 53.280 57.040 54.180 57.940 ;
        RECT 63.720 56.780 64.940 57.440 ;
        RECT 69.760 56.800 70.980 57.460 ;
        RECT 71.640 56.800 72.860 57.460 ;
        RECT 73.520 56.810 74.740 57.470 ;
        RECT 75.940 57.040 76.840 57.940 ;
        RECT 86.380 56.780 87.600 57.440 ;
        RECT 92.420 56.800 93.640 57.460 ;
        RECT 94.300 56.800 95.520 57.460 ;
        RECT 96.180 56.810 97.400 57.470 ;
        RECT 98.600 57.040 99.500 57.940 ;
        RECT 109.040 56.780 110.260 57.440 ;
        RECT 115.080 56.800 116.300 57.460 ;
        RECT 116.960 56.800 118.180 57.460 ;
        RECT 118.840 56.810 120.060 57.470 ;
        RECT 121.260 57.040 122.160 57.940 ;
        RECT 30.945 54.445 31.895 55.395 ;
        RECT 127.800 54.430 128.800 55.430 ;
      LAYER met3 ;
        RECT 59.500 183.705 61.080 184.035 ;
        RECT 78.010 183.705 79.590 184.035 ;
        RECT 96.520 183.705 98.100 184.035 ;
        RECT 115.030 183.705 116.610 184.035 ;
        RECT 59.500 178.265 61.080 178.595 ;
        RECT 78.010 178.265 79.590 178.595 ;
        RECT 96.520 178.265 98.100 178.595 ;
        RECT 115.030 178.265 116.610 178.595 ;
        RECT 59.500 172.825 61.080 173.155 ;
        RECT 78.010 172.825 79.590 173.155 ;
        RECT 96.520 172.825 98.100 173.155 ;
        RECT 115.030 172.825 116.610 173.155 ;
        RECT 59.500 167.385 61.080 167.715 ;
        RECT 78.010 167.385 79.590 167.715 ;
        RECT 96.520 167.385 98.100 167.715 ;
        RECT 115.030 167.385 116.610 167.715 ;
        RECT 59.500 161.945 61.080 162.275 ;
        RECT 78.010 161.945 79.590 162.275 ;
        RECT 96.520 161.945 98.100 162.275 ;
        RECT 115.030 161.945 116.610 162.275 ;
        RECT 59.500 156.505 61.080 156.835 ;
        RECT 78.010 156.505 79.590 156.835 ;
        RECT 96.520 156.505 98.100 156.835 ;
        RECT 115.030 156.505 116.610 156.835 ;
        RECT 12.000 147.000 116.620 148.600 ;
        RECT 63.830 127.510 64.830 127.630 ;
        RECT 69.870 127.530 70.870 127.650 ;
        RECT 71.750 127.530 72.750 127.650 ;
        RECT 73.630 127.540 74.630 127.660 ;
        RECT 63.670 126.750 64.990 127.510 ;
        RECT 69.710 126.770 71.030 127.530 ;
        RECT 71.590 126.770 72.910 127.530 ;
        RECT 73.470 126.780 74.790 127.540 ;
        RECT 30.895 125.440 31.945 125.455 ;
        RECT 63.830 125.440 64.830 126.750 ;
        RECT 69.870 125.440 70.870 126.770 ;
        RECT 71.750 125.440 72.750 126.770 ;
        RECT 73.630 125.440 74.630 126.780 ;
        RECT 75.890 125.440 76.890 128.010 ;
        RECT 86.490 127.510 87.490 127.630 ;
        RECT 92.530 127.530 93.530 127.650 ;
        RECT 94.410 127.530 95.410 127.650 ;
        RECT 96.290 127.540 97.290 127.660 ;
        RECT 86.330 126.750 87.650 127.510 ;
        RECT 92.370 126.770 93.690 127.530 ;
        RECT 94.250 126.770 95.570 127.530 ;
        RECT 96.130 126.780 97.450 127.540 ;
        RECT 86.490 125.440 87.490 126.750 ;
        RECT 92.530 125.440 93.530 126.770 ;
        RECT 94.410 125.440 95.410 126.770 ;
        RECT 96.290 125.440 97.290 126.780 ;
        RECT 98.550 125.440 99.550 128.010 ;
        RECT 109.150 127.510 110.150 127.630 ;
        RECT 115.190 127.530 116.190 127.650 ;
        RECT 117.070 127.530 118.070 127.650 ;
        RECT 118.950 127.540 119.950 127.660 ;
        RECT 108.990 126.750 110.310 127.510 ;
        RECT 115.030 126.770 116.350 127.530 ;
        RECT 116.910 126.770 118.230 127.530 ;
        RECT 118.790 126.780 120.110 127.540 ;
        RECT 109.150 125.440 110.150 126.750 ;
        RECT 115.190 125.440 116.190 126.770 ;
        RECT 117.070 125.440 118.070 126.770 ;
        RECT 118.950 125.440 119.950 126.780 ;
        RECT 121.210 125.440 122.210 128.010 ;
        RECT 123.875 125.440 124.875 128.810 ;
        RECT 127.775 125.440 128.825 125.465 ;
        RECT 30.870 124.440 128.830 125.440 ;
        RECT 30.895 124.405 31.945 124.440 ;
        RECT 61.250 121.580 62.250 124.440 ;
        RECT 83.910 121.580 84.910 124.440 ;
        RECT 106.570 121.580 107.570 124.440 ;
        RECT 127.775 124.415 128.825 124.440 ;
        RECT 41.170 110.170 42.170 110.290 ;
        RECT 47.210 110.190 48.210 110.310 ;
        RECT 49.090 110.190 50.090 110.310 ;
        RECT 50.970 110.200 51.970 110.320 ;
        RECT 41.010 109.410 42.330 110.170 ;
        RECT 47.050 109.430 48.370 110.190 ;
        RECT 48.930 109.430 50.250 110.190 ;
        RECT 50.810 109.440 52.130 110.200 ;
        RECT 30.895 108.100 31.945 108.145 ;
        RECT 41.170 108.100 42.170 109.410 ;
        RECT 47.210 108.100 48.210 109.430 ;
        RECT 49.090 108.100 50.090 109.430 ;
        RECT 50.970 108.100 51.970 109.440 ;
        RECT 53.230 108.100 54.230 110.670 ;
        RECT 63.830 110.170 64.830 110.290 ;
        RECT 69.870 110.190 70.870 110.310 ;
        RECT 71.750 110.190 72.750 110.310 ;
        RECT 73.630 110.200 74.630 110.320 ;
        RECT 63.670 109.410 64.990 110.170 ;
        RECT 69.710 109.430 71.030 110.190 ;
        RECT 71.590 109.430 72.910 110.190 ;
        RECT 73.470 109.440 74.790 110.200 ;
        RECT 63.830 108.100 64.830 109.410 ;
        RECT 69.870 108.100 70.870 109.430 ;
        RECT 71.750 108.100 72.750 109.430 ;
        RECT 73.630 108.100 74.630 109.440 ;
        RECT 75.890 108.100 76.890 110.670 ;
        RECT 86.490 110.170 87.490 110.290 ;
        RECT 92.530 110.190 93.530 110.310 ;
        RECT 94.410 110.190 95.410 110.310 ;
        RECT 96.290 110.200 97.290 110.320 ;
        RECT 86.330 109.410 87.650 110.170 ;
        RECT 92.370 109.430 93.690 110.190 ;
        RECT 94.250 109.430 95.570 110.190 ;
        RECT 96.130 109.440 97.450 110.200 ;
        RECT 86.490 108.100 87.490 109.410 ;
        RECT 92.530 108.100 93.530 109.430 ;
        RECT 94.410 108.100 95.410 109.430 ;
        RECT 96.290 108.100 97.290 109.440 ;
        RECT 98.550 108.100 99.550 110.670 ;
        RECT 109.150 110.170 110.150 110.290 ;
        RECT 115.190 110.190 116.190 110.310 ;
        RECT 117.070 110.190 118.070 110.310 ;
        RECT 118.950 110.200 119.950 110.320 ;
        RECT 108.990 109.410 110.310 110.170 ;
        RECT 115.030 109.430 116.350 110.190 ;
        RECT 116.910 109.430 118.230 110.190 ;
        RECT 118.790 109.440 120.110 110.200 ;
        RECT 109.150 108.100 110.150 109.410 ;
        RECT 115.190 108.100 116.190 109.430 ;
        RECT 117.070 108.100 118.070 109.430 ;
        RECT 118.950 108.100 119.950 109.440 ;
        RECT 121.210 108.100 122.210 110.670 ;
        RECT 127.775 108.100 128.825 108.125 ;
        RECT 30.870 107.100 128.830 108.100 ;
        RECT 30.895 107.095 31.945 107.100 ;
        RECT 38.590 104.240 39.590 107.100 ;
        RECT 61.250 104.240 62.250 107.100 ;
        RECT 83.910 104.240 84.910 107.100 ;
        RECT 106.570 104.240 107.570 107.100 ;
        RECT 127.775 107.075 128.825 107.100 ;
        RECT 41.170 92.830 42.170 92.950 ;
        RECT 47.210 92.850 48.210 92.970 ;
        RECT 49.090 92.850 50.090 92.970 ;
        RECT 50.970 92.860 51.970 92.980 ;
        RECT 41.010 92.070 42.330 92.830 ;
        RECT 47.050 92.090 48.370 92.850 ;
        RECT 48.930 92.090 50.250 92.850 ;
        RECT 50.810 92.100 52.130 92.860 ;
        RECT 30.895 90.760 31.945 90.785 ;
        RECT 41.170 90.760 42.170 92.070 ;
        RECT 47.210 90.760 48.210 92.090 ;
        RECT 49.090 90.760 50.090 92.090 ;
        RECT 50.970 90.760 51.970 92.100 ;
        RECT 53.230 90.760 54.230 93.330 ;
        RECT 63.830 92.830 64.830 92.950 ;
        RECT 69.870 92.850 70.870 92.970 ;
        RECT 71.750 92.850 72.750 92.970 ;
        RECT 73.630 92.860 74.630 92.980 ;
        RECT 63.670 92.070 64.990 92.830 ;
        RECT 69.710 92.090 71.030 92.850 ;
        RECT 71.590 92.090 72.910 92.850 ;
        RECT 73.470 92.100 74.790 92.860 ;
        RECT 63.830 90.760 64.830 92.070 ;
        RECT 69.870 90.760 70.870 92.090 ;
        RECT 71.750 90.760 72.750 92.090 ;
        RECT 73.630 90.760 74.630 92.100 ;
        RECT 75.890 90.760 76.890 93.330 ;
        RECT 86.490 92.830 87.490 92.950 ;
        RECT 92.530 92.850 93.530 92.970 ;
        RECT 94.410 92.850 95.410 92.970 ;
        RECT 96.290 92.860 97.290 92.980 ;
        RECT 86.330 92.070 87.650 92.830 ;
        RECT 92.370 92.090 93.690 92.850 ;
        RECT 94.250 92.090 95.570 92.850 ;
        RECT 96.130 92.100 97.450 92.860 ;
        RECT 86.490 90.760 87.490 92.070 ;
        RECT 92.530 90.760 93.530 92.090 ;
        RECT 94.410 90.760 95.410 92.090 ;
        RECT 96.290 90.760 97.290 92.100 ;
        RECT 98.550 90.760 99.550 93.330 ;
        RECT 109.150 92.830 110.150 92.950 ;
        RECT 115.190 92.850 116.190 92.970 ;
        RECT 117.070 92.850 118.070 92.970 ;
        RECT 118.950 92.860 119.950 92.980 ;
        RECT 108.990 92.070 110.310 92.830 ;
        RECT 115.030 92.090 116.350 92.850 ;
        RECT 116.910 92.090 118.230 92.850 ;
        RECT 118.790 92.100 120.110 92.860 ;
        RECT 109.150 90.760 110.150 92.070 ;
        RECT 115.190 90.760 116.190 92.090 ;
        RECT 117.070 90.760 118.070 92.090 ;
        RECT 118.950 90.760 119.950 92.100 ;
        RECT 121.210 90.760 122.210 93.330 ;
        RECT 127.775 90.760 128.825 90.775 ;
        RECT 30.870 89.760 128.830 90.760 ;
        RECT 30.895 89.735 31.945 89.760 ;
        RECT 38.590 86.900 39.590 89.760 ;
        RECT 61.250 86.900 62.250 89.760 ;
        RECT 83.910 86.900 84.910 89.760 ;
        RECT 106.570 86.900 107.570 89.760 ;
        RECT 127.775 89.725 128.825 89.760 ;
        RECT 41.170 75.490 42.170 75.610 ;
        RECT 47.210 75.510 48.210 75.630 ;
        RECT 49.090 75.510 50.090 75.630 ;
        RECT 50.970 75.520 51.970 75.640 ;
        RECT 41.010 74.730 42.330 75.490 ;
        RECT 47.050 74.750 48.370 75.510 ;
        RECT 48.930 74.750 50.250 75.510 ;
        RECT 50.810 74.760 52.130 75.520 ;
        RECT 30.895 73.420 31.945 73.465 ;
        RECT 41.170 73.420 42.170 74.730 ;
        RECT 47.210 73.420 48.210 74.750 ;
        RECT 49.090 73.420 50.090 74.750 ;
        RECT 50.970 73.420 51.970 74.760 ;
        RECT 53.230 73.420 54.230 75.990 ;
        RECT 63.830 75.490 64.830 75.610 ;
        RECT 69.870 75.510 70.870 75.630 ;
        RECT 71.750 75.510 72.750 75.630 ;
        RECT 73.630 75.520 74.630 75.640 ;
        RECT 63.670 74.730 64.990 75.490 ;
        RECT 69.710 74.750 71.030 75.510 ;
        RECT 71.590 74.750 72.910 75.510 ;
        RECT 73.470 74.760 74.790 75.520 ;
        RECT 63.830 73.420 64.830 74.730 ;
        RECT 69.870 73.420 70.870 74.750 ;
        RECT 71.750 73.420 72.750 74.750 ;
        RECT 73.630 73.420 74.630 74.760 ;
        RECT 75.890 73.420 76.890 75.990 ;
        RECT 86.490 75.490 87.490 75.610 ;
        RECT 92.530 75.510 93.530 75.630 ;
        RECT 94.410 75.510 95.410 75.630 ;
        RECT 96.290 75.520 97.290 75.640 ;
        RECT 86.330 74.730 87.650 75.490 ;
        RECT 92.370 74.750 93.690 75.510 ;
        RECT 94.250 74.750 95.570 75.510 ;
        RECT 96.130 74.760 97.450 75.520 ;
        RECT 86.490 73.420 87.490 74.730 ;
        RECT 92.530 73.420 93.530 74.750 ;
        RECT 94.410 73.420 95.410 74.750 ;
        RECT 96.290 73.420 97.290 74.760 ;
        RECT 98.550 73.420 99.550 75.990 ;
        RECT 109.150 75.490 110.150 75.610 ;
        RECT 115.190 75.510 116.190 75.630 ;
        RECT 117.070 75.510 118.070 75.630 ;
        RECT 118.950 75.520 119.950 75.640 ;
        RECT 108.990 74.730 110.310 75.490 ;
        RECT 115.030 74.750 116.350 75.510 ;
        RECT 116.910 74.750 118.230 75.510 ;
        RECT 118.790 74.760 120.110 75.520 ;
        RECT 109.150 73.420 110.150 74.730 ;
        RECT 115.190 73.420 116.190 74.750 ;
        RECT 117.070 73.420 118.070 74.750 ;
        RECT 118.950 73.420 119.950 74.760 ;
        RECT 121.210 73.420 122.210 75.990 ;
        RECT 127.775 73.420 128.825 73.445 ;
        RECT 30.870 72.420 128.830 73.420 ;
        RECT 30.895 72.415 31.945 72.420 ;
        RECT 38.590 69.560 39.590 72.420 ;
        RECT 61.250 69.560 62.250 72.420 ;
        RECT 83.910 69.560 84.910 72.420 ;
        RECT 106.570 69.560 107.570 72.420 ;
        RECT 127.775 72.395 128.825 72.420 ;
        RECT 41.170 57.490 42.170 57.610 ;
        RECT 47.210 57.510 48.210 57.630 ;
        RECT 49.090 57.510 50.090 57.630 ;
        RECT 50.970 57.520 51.970 57.640 ;
        RECT 41.010 56.730 42.330 57.490 ;
        RECT 47.050 56.750 48.370 57.510 ;
        RECT 48.930 56.750 50.250 57.510 ;
        RECT 50.810 56.760 52.130 57.520 ;
        RECT 41.170 55.420 42.170 56.730 ;
        RECT 47.210 55.420 48.210 56.750 ;
        RECT 49.090 55.420 50.090 56.750 ;
        RECT 50.970 55.420 51.970 56.760 ;
        RECT 53.230 55.420 54.230 57.990 ;
        RECT 63.830 57.490 64.830 57.610 ;
        RECT 69.870 57.510 70.870 57.630 ;
        RECT 71.750 57.510 72.750 57.630 ;
        RECT 73.630 57.520 74.630 57.640 ;
        RECT 63.670 56.730 64.990 57.490 ;
        RECT 69.710 56.750 71.030 57.510 ;
        RECT 71.590 56.750 72.910 57.510 ;
        RECT 73.470 56.760 74.790 57.520 ;
        RECT 63.830 55.420 64.830 56.730 ;
        RECT 69.870 55.420 70.870 56.750 ;
        RECT 71.750 55.420 72.750 56.750 ;
        RECT 73.630 55.420 74.630 56.760 ;
        RECT 75.890 55.420 76.890 57.990 ;
        RECT 86.490 57.490 87.490 57.610 ;
        RECT 92.530 57.510 93.530 57.630 ;
        RECT 94.410 57.510 95.410 57.630 ;
        RECT 96.290 57.520 97.290 57.640 ;
        RECT 86.330 56.730 87.650 57.490 ;
        RECT 92.370 56.750 93.690 57.510 ;
        RECT 94.250 56.750 95.570 57.510 ;
        RECT 96.130 56.760 97.450 57.520 ;
        RECT 86.490 55.420 87.490 56.730 ;
        RECT 92.530 55.420 93.530 56.750 ;
        RECT 94.410 55.420 95.410 56.750 ;
        RECT 96.290 55.420 97.290 56.760 ;
        RECT 98.550 55.420 99.550 57.990 ;
        RECT 109.150 57.490 110.150 57.610 ;
        RECT 115.190 57.510 116.190 57.630 ;
        RECT 117.070 57.510 118.070 57.630 ;
        RECT 118.950 57.520 119.950 57.640 ;
        RECT 108.990 56.730 110.310 57.490 ;
        RECT 115.030 56.750 116.350 57.510 ;
        RECT 116.910 56.750 118.230 57.510 ;
        RECT 118.790 56.760 120.110 57.520 ;
        RECT 109.150 55.420 110.150 56.730 ;
        RECT 115.190 55.420 116.190 56.750 ;
        RECT 117.070 55.420 118.070 56.750 ;
        RECT 118.950 55.420 119.950 56.760 ;
        RECT 121.210 55.420 122.210 57.990 ;
        RECT 127.775 55.420 128.825 55.455 ;
        RECT 30.870 54.420 128.830 55.420 ;
        RECT 127.775 54.405 128.825 54.420 ;
      LAYER via3 ;
        RECT 59.530 183.710 59.850 184.030 ;
        RECT 59.930 183.710 60.250 184.030 ;
        RECT 60.330 183.710 60.650 184.030 ;
        RECT 60.730 183.710 61.050 184.030 ;
        RECT 78.040 183.710 78.360 184.030 ;
        RECT 78.440 183.710 78.760 184.030 ;
        RECT 78.840 183.710 79.160 184.030 ;
        RECT 79.240 183.710 79.560 184.030 ;
        RECT 96.550 183.710 96.870 184.030 ;
        RECT 96.950 183.710 97.270 184.030 ;
        RECT 97.350 183.710 97.670 184.030 ;
        RECT 97.750 183.710 98.070 184.030 ;
        RECT 115.060 183.710 115.380 184.030 ;
        RECT 115.460 183.710 115.780 184.030 ;
        RECT 115.860 183.710 116.180 184.030 ;
        RECT 116.260 183.710 116.580 184.030 ;
        RECT 59.530 178.270 59.850 178.590 ;
        RECT 59.930 178.270 60.250 178.590 ;
        RECT 60.330 178.270 60.650 178.590 ;
        RECT 60.730 178.270 61.050 178.590 ;
        RECT 78.040 178.270 78.360 178.590 ;
        RECT 78.440 178.270 78.760 178.590 ;
        RECT 78.840 178.270 79.160 178.590 ;
        RECT 79.240 178.270 79.560 178.590 ;
        RECT 96.550 178.270 96.870 178.590 ;
        RECT 96.950 178.270 97.270 178.590 ;
        RECT 97.350 178.270 97.670 178.590 ;
        RECT 97.750 178.270 98.070 178.590 ;
        RECT 115.060 178.270 115.380 178.590 ;
        RECT 115.460 178.270 115.780 178.590 ;
        RECT 115.860 178.270 116.180 178.590 ;
        RECT 116.260 178.270 116.580 178.590 ;
        RECT 59.530 172.830 59.850 173.150 ;
        RECT 59.930 172.830 60.250 173.150 ;
        RECT 60.330 172.830 60.650 173.150 ;
        RECT 60.730 172.830 61.050 173.150 ;
        RECT 78.040 172.830 78.360 173.150 ;
        RECT 78.440 172.830 78.760 173.150 ;
        RECT 78.840 172.830 79.160 173.150 ;
        RECT 79.240 172.830 79.560 173.150 ;
        RECT 96.550 172.830 96.870 173.150 ;
        RECT 96.950 172.830 97.270 173.150 ;
        RECT 97.350 172.830 97.670 173.150 ;
        RECT 97.750 172.830 98.070 173.150 ;
        RECT 115.060 172.830 115.380 173.150 ;
        RECT 115.460 172.830 115.780 173.150 ;
        RECT 115.860 172.830 116.180 173.150 ;
        RECT 116.260 172.830 116.580 173.150 ;
        RECT 59.530 167.390 59.850 167.710 ;
        RECT 59.930 167.390 60.250 167.710 ;
        RECT 60.330 167.390 60.650 167.710 ;
        RECT 60.730 167.390 61.050 167.710 ;
        RECT 78.040 167.390 78.360 167.710 ;
        RECT 78.440 167.390 78.760 167.710 ;
        RECT 78.840 167.390 79.160 167.710 ;
        RECT 79.240 167.390 79.560 167.710 ;
        RECT 96.550 167.390 96.870 167.710 ;
        RECT 96.950 167.390 97.270 167.710 ;
        RECT 97.350 167.390 97.670 167.710 ;
        RECT 97.750 167.390 98.070 167.710 ;
        RECT 115.060 167.390 115.380 167.710 ;
        RECT 115.460 167.390 115.780 167.710 ;
        RECT 115.860 167.390 116.180 167.710 ;
        RECT 116.260 167.390 116.580 167.710 ;
        RECT 59.530 161.950 59.850 162.270 ;
        RECT 59.930 161.950 60.250 162.270 ;
        RECT 60.330 161.950 60.650 162.270 ;
        RECT 60.730 161.950 61.050 162.270 ;
        RECT 78.040 161.950 78.360 162.270 ;
        RECT 78.440 161.950 78.760 162.270 ;
        RECT 78.840 161.950 79.160 162.270 ;
        RECT 79.240 161.950 79.560 162.270 ;
        RECT 96.550 161.950 96.870 162.270 ;
        RECT 96.950 161.950 97.270 162.270 ;
        RECT 97.350 161.950 97.670 162.270 ;
        RECT 97.750 161.950 98.070 162.270 ;
        RECT 115.060 161.950 115.380 162.270 ;
        RECT 115.460 161.950 115.780 162.270 ;
        RECT 115.860 161.950 116.180 162.270 ;
        RECT 116.260 161.950 116.580 162.270 ;
        RECT 59.530 156.510 59.850 156.830 ;
        RECT 59.930 156.510 60.250 156.830 ;
        RECT 60.330 156.510 60.650 156.830 ;
        RECT 60.730 156.510 61.050 156.830 ;
        RECT 78.040 156.510 78.360 156.830 ;
        RECT 78.440 156.510 78.760 156.830 ;
        RECT 78.840 156.510 79.160 156.830 ;
        RECT 79.240 156.510 79.560 156.830 ;
        RECT 96.550 156.510 96.870 156.830 ;
        RECT 96.950 156.510 97.270 156.830 ;
        RECT 97.350 156.510 97.670 156.830 ;
        RECT 97.750 156.510 98.070 156.830 ;
        RECT 115.060 156.510 115.380 156.830 ;
        RECT 115.460 156.510 115.780 156.830 ;
        RECT 115.860 156.510 116.180 156.830 ;
        RECT 116.260 156.510 116.580 156.830 ;
        RECT 22.100 147.100 23.500 148.500 ;
        RECT 59.595 147.100 60.995 148.500 ;
        RECT 78.105 147.100 79.505 148.500 ;
        RECT 96.615 147.100 98.015 148.500 ;
        RECT 115.125 147.100 116.525 148.500 ;
        RECT 59.590 124.540 60.990 125.350 ;
        RECT 78.100 124.540 79.500 125.350 ;
        RECT 96.610 124.540 98.010 125.350 ;
        RECT 115.120 124.540 116.520 125.350 ;
        RECT 59.590 107.200 60.990 108.010 ;
        RECT 78.100 107.200 79.500 108.010 ;
        RECT 96.610 107.200 98.010 108.010 ;
        RECT 115.120 107.200 116.520 108.010 ;
        RECT 59.590 89.860 60.990 90.670 ;
        RECT 78.100 89.860 79.500 90.670 ;
        RECT 96.610 89.860 98.010 90.670 ;
        RECT 115.120 89.860 116.520 90.670 ;
        RECT 59.590 72.520 60.990 73.330 ;
        RECT 78.100 72.520 79.500 73.330 ;
        RECT 96.610 72.520 98.010 73.330 ;
        RECT 115.120 72.520 116.520 73.330 ;
        RECT 59.590 54.520 60.990 55.330 ;
        RECT 78.100 54.520 79.500 55.330 ;
        RECT 96.610 54.520 98.010 55.330 ;
        RECT 115.120 54.520 116.520 55.330 ;
      LAYER met4 ;
        RECT 22.000 5.000 23.600 220.760 ;
        RECT 59.490 44.400 61.090 186.850 ;
        RECT 78.000 44.400 79.600 186.850 ;
        RECT 96.510 44.400 98.110 186.850 ;
        RECT 115.020 44.400 116.620 186.850 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 41.785 183.975 43.155 184.785 ;
        RECT 48.250 184.655 49.595 184.885 ;
        RECT 50.550 184.655 51.895 184.885 ;
        RECT 52.390 184.655 53.735 184.885 ;
        RECT 44.085 183.975 46.825 184.655 ;
        RECT 47.765 183.975 49.595 184.655 ;
        RECT 50.065 183.975 51.895 184.655 ;
        RECT 51.905 183.975 53.735 184.655 ;
        RECT 55.125 184.655 56.470 184.885 ;
        RECT 57.910 184.655 59.255 184.885 ;
        RECT 59.750 184.655 61.095 184.885 ;
        RECT 55.125 183.975 56.955 184.655 ;
        RECT 57.425 183.975 59.255 184.655 ;
        RECT 59.265 183.975 61.095 184.655 ;
        RECT 61.105 184.655 62.450 184.885 ;
        RECT 66.190 184.655 67.535 184.885 ;
        RECT 61.105 183.975 62.935 184.655 ;
        RECT 62.945 183.975 65.685 184.655 ;
        RECT 65.705 183.975 67.535 184.655 ;
        RECT 68.005 184.655 69.350 184.885 ;
        RECT 70.330 184.655 71.675 184.885 ;
        RECT 68.005 183.975 69.835 184.655 ;
        RECT 69.845 183.975 71.675 184.655 ;
        RECT 71.685 184.655 73.030 184.885 ;
        RECT 74.445 184.655 75.790 184.885 ;
        RECT 76.745 184.655 78.090 184.885 ;
        RECT 71.685 183.975 73.515 184.655 ;
        RECT 74.445 183.975 76.275 184.655 ;
        RECT 76.745 183.975 78.575 184.655 ;
        RECT 78.585 183.975 80.415 184.785 ;
        RECT 81.945 183.975 84.555 184.885 ;
        RECT 84.575 183.975 87.315 184.655 ;
        RECT 87.325 183.975 88.695 184.755 ;
        RECT 89.165 183.975 90.535 184.755 ;
        RECT 91.005 183.975 92.375 184.755 ;
        RECT 93.765 183.975 97.635 184.885 ;
        RECT 104.785 184.655 105.715 184.885 ;
        RECT 98.835 183.975 101.575 184.655 ;
        RECT 101.815 183.975 105.715 184.655 ;
        RECT 107.565 184.655 108.910 184.885 ;
        RECT 109.405 184.655 110.335 184.885 ;
        RECT 107.565 183.975 109.395 184.655 ;
        RECT 109.405 183.975 113.305 184.655 ;
        RECT 114.465 183.975 115.835 184.785 ;
        RECT 41.925 183.765 42.095 183.975 ;
        RECT 43.315 183.810 43.475 183.930 ;
        RECT 44.225 183.785 44.395 183.975 ;
        RECT 45.605 183.765 45.775 183.955 ;
        RECT 46.065 183.765 46.235 183.955 ;
        RECT 46.995 183.820 47.155 183.930 ;
        RECT 47.905 183.765 48.075 183.975 ;
        RECT 49.740 183.815 49.860 183.925 ;
        RECT 50.205 183.785 50.375 183.975 ;
        RECT 52.045 183.785 52.215 183.975 ;
        RECT 41.785 182.955 43.155 183.765 ;
        RECT 44.085 183.085 45.915 183.765 ;
        RECT 45.925 183.085 47.755 183.765 ;
        RECT 44.085 182.855 45.430 183.085 ;
        RECT 46.410 182.855 47.755 183.085 ;
        RECT 47.765 182.955 53.275 183.765 ;
        RECT 53.430 183.735 53.600 183.955 ;
        RECT 53.895 183.820 54.055 183.930 ;
        RECT 56.645 183.785 56.815 183.975 ;
        RECT 57.100 183.815 57.220 183.925 ;
        RECT 57.565 183.785 57.735 183.975 ;
        RECT 59.405 183.955 59.575 183.975 ;
        RECT 59.400 183.785 59.575 183.955 ;
        RECT 59.400 183.765 59.570 183.785 ;
        RECT 59.865 183.765 60.035 183.955 ;
        RECT 62.625 183.785 62.795 183.975 ;
        RECT 63.085 183.785 63.255 183.975 ;
        RECT 65.845 183.785 66.015 183.975 ;
        RECT 66.950 183.765 67.120 183.955 ;
        RECT 68.155 183.810 68.315 183.920 ;
        RECT 69.525 183.785 69.695 183.975 ;
        RECT 69.985 183.785 70.155 183.975 ;
        RECT 72.470 183.765 72.640 183.955 ;
        RECT 73.205 183.785 73.375 183.975 ;
        RECT 73.675 183.820 73.835 183.930 ;
        RECT 75.965 183.785 76.135 183.975 ;
        RECT 76.420 183.815 76.540 183.925 ;
        RECT 76.610 183.765 76.780 183.955 ;
        RECT 78.265 183.785 78.435 183.975 ;
        RECT 78.725 183.785 78.895 183.975 ;
        RECT 81.035 183.820 81.195 183.930 ;
        RECT 81.510 183.785 81.680 183.955 ;
        RECT 81.510 183.765 81.620 183.785 ;
        RECT 82.220 183.765 82.390 183.955 ;
        RECT 84.240 183.785 84.410 183.975 ;
        RECT 86.085 183.765 86.255 183.955 ;
        RECT 87.005 183.785 87.175 183.975 ;
        RECT 88.200 183.765 88.370 183.955 ;
        RECT 88.375 183.785 88.545 183.975 ;
        RECT 88.840 183.815 88.960 183.925 ;
        RECT 90.225 183.785 90.395 183.975 ;
        RECT 90.680 183.815 90.800 183.925 ;
        RECT 92.055 183.785 92.225 183.975 ;
        RECT 97.580 183.955 97.635 183.975 ;
        RECT 92.535 183.820 92.695 183.930 ;
        RECT 92.985 183.765 93.155 183.955 ;
        RECT 94.180 183.765 94.350 183.955 ;
        RECT 97.580 183.785 97.750 183.955 ;
        RECT 98.055 183.820 98.215 183.930 ;
        RECT 98.320 183.765 98.490 183.955 ;
        RECT 101.265 183.785 101.435 183.975 ;
        RECT 102.180 183.815 102.300 183.925 ;
        RECT 105.130 183.785 105.300 183.975 ;
        RECT 105.860 183.815 105.980 183.925 ;
        RECT 106.320 183.785 106.490 183.955 ;
        RECT 106.795 183.820 106.955 183.930 ;
        RECT 106.320 183.765 106.375 183.785 ;
        RECT 107.060 183.765 107.230 183.955 ;
        RECT 109.085 183.785 109.255 183.975 ;
        RECT 109.820 183.785 109.990 183.975 ;
        RECT 110.930 183.765 111.100 183.955 ;
        RECT 113.695 183.810 113.855 183.930 ;
        RECT 115.525 183.765 115.695 183.975 ;
        RECT 55.560 183.735 56.495 183.765 ;
        RECT 53.430 183.535 56.495 183.735 ;
        RECT 53.285 183.055 56.495 183.535 ;
        RECT 53.285 182.855 54.215 183.055 ;
        RECT 55.545 182.855 56.495 183.055 ;
        RECT 56.505 182.855 59.715 183.765 ;
        RECT 59.725 182.955 63.395 183.765 ;
        RECT 63.635 183.085 67.535 183.765 ;
        RECT 69.155 183.085 73.055 183.765 ;
        RECT 73.295 183.085 77.195 183.765 ;
        RECT 66.605 182.855 67.535 183.085 ;
        RECT 72.125 182.855 73.055 183.085 ;
        RECT 76.265 182.855 77.195 183.085 ;
        RECT 77.205 183.085 81.620 183.765 ;
        RECT 81.805 183.085 85.705 183.765 ;
        RECT 77.205 182.855 81.135 183.085 ;
        RECT 81.805 182.855 82.735 183.085 ;
        RECT 85.945 182.955 87.775 183.765 ;
        RECT 87.785 183.085 91.685 183.765 ;
        RECT 87.785 182.855 88.715 183.085 ;
        RECT 91.925 182.985 93.295 183.765 ;
        RECT 93.765 183.085 97.665 183.765 ;
        RECT 97.905 183.085 101.805 183.765 ;
        RECT 93.765 182.855 94.695 183.085 ;
        RECT 97.905 182.855 98.835 183.085 ;
        RECT 102.505 182.855 106.375 183.765 ;
        RECT 106.645 183.085 110.545 183.765 ;
        RECT 106.645 182.855 107.575 183.085 ;
        RECT 110.785 182.855 113.395 183.765 ;
        RECT 114.465 182.955 115.835 183.765 ;
        RECT 41.785 178.535 43.155 179.345 ;
        RECT 43.165 178.535 48.675 179.345 ;
        RECT 49.685 178.535 53.135 179.445 ;
        RECT 53.295 178.535 54.645 179.445 ;
        RECT 55.125 178.535 60.635 179.345 ;
        RECT 60.645 178.535 62.475 179.345 ;
        RECT 62.945 179.215 63.875 179.445 ;
        RECT 62.945 178.535 66.845 179.215 ;
        RECT 68.005 178.535 69.375 179.315 ;
        RECT 69.385 178.535 70.755 179.345 ;
        RECT 70.815 178.535 73.005 179.445 ;
        RECT 73.065 178.535 74.895 179.345 ;
        RECT 74.905 178.535 76.735 179.215 ;
        RECT 76.745 178.535 80.415 179.345 ;
        RECT 80.885 178.535 86.395 179.345 ;
        RECT 86.405 178.535 88.235 179.345 ;
        RECT 91.905 179.215 92.835 179.445 ;
        RECT 88.935 178.535 92.835 179.215 ;
        RECT 92.845 178.535 94.215 179.315 ;
        RECT 95.145 179.215 96.490 179.445 ;
        RECT 95.145 178.535 96.975 179.215 ;
        RECT 96.985 178.535 98.355 179.315 ;
        RECT 98.365 178.535 99.735 179.315 ;
        RECT 100.205 179.215 101.135 179.445 ;
        RECT 100.205 178.535 104.105 179.215 ;
        RECT 104.345 178.535 105.715 179.315 ;
        RECT 109.605 179.215 113.535 179.445 ;
        RECT 106.645 178.535 108.475 179.215 ;
        RECT 109.120 178.535 113.535 179.215 ;
        RECT 114.465 178.535 115.835 179.345 ;
        RECT 41.925 178.325 42.095 178.535 ;
        RECT 43.305 178.325 43.475 178.535 ;
        RECT 48.835 178.370 48.995 178.490 ;
        RECT 49.745 178.325 49.915 178.535 ;
        RECT 52.505 178.325 52.675 178.515 ;
        RECT 54.345 178.345 54.515 178.535 ;
        RECT 55.265 178.345 55.435 178.535 ;
        RECT 58.020 178.375 58.140 178.485 ;
        RECT 58.760 178.325 58.930 178.515 ;
        RECT 60.785 178.345 60.955 178.535 ;
        RECT 62.625 178.485 62.795 178.515 ;
        RECT 62.620 178.375 62.795 178.485 ;
        RECT 62.625 178.325 62.795 178.375 ;
        RECT 63.360 178.345 63.530 178.535 ;
        RECT 65.385 178.325 65.555 178.515 ;
        RECT 67.235 178.485 67.395 178.490 ;
        RECT 67.220 178.380 67.395 178.485 ;
        RECT 67.220 178.375 67.340 178.380 ;
        RECT 69.055 178.345 69.225 178.535 ;
        RECT 69.525 178.345 69.695 178.535 ;
        RECT 69.980 178.325 70.150 178.515 ;
        RECT 70.445 178.325 70.615 178.515 ;
        RECT 72.745 178.345 72.915 178.535 ;
        RECT 73.205 178.345 73.375 178.535 ;
        RECT 76.240 178.325 76.410 178.515 ;
        RECT 76.425 178.345 76.595 178.535 ;
        RECT 76.885 178.345 77.055 178.535 ;
        RECT 81.025 178.345 81.195 178.535 ;
        RECT 86.545 178.345 86.715 178.535 ;
        RECT 88.380 178.375 88.500 178.485 ;
        RECT 89.305 178.325 89.475 178.515 ;
        RECT 91.605 178.345 91.775 178.515 ;
        RECT 91.605 178.325 91.755 178.345 ;
        RECT 92.065 178.325 92.235 178.515 ;
        RECT 92.250 178.345 92.420 178.535 ;
        RECT 92.995 178.345 93.165 178.535 ;
        RECT 94.180 178.325 94.350 178.515 ;
        RECT 94.375 178.380 94.535 178.490 ;
        RECT 96.665 178.345 96.835 178.535 ;
        RECT 98.045 178.515 98.215 178.535 ;
        RECT 98.045 178.345 98.220 178.515 ;
        RECT 99.425 178.345 99.595 178.535 ;
        RECT 99.880 178.375 100.000 178.485 ;
        RECT 100.620 178.345 100.790 178.535 ;
        RECT 102.195 178.370 102.355 178.480 ;
        RECT 98.165 178.325 98.220 178.345 ;
        RECT 103.380 178.325 103.550 178.515 ;
        RECT 105.395 178.345 105.565 178.535 ;
        RECT 105.860 178.375 105.980 178.485 ;
        RECT 106.785 178.345 106.955 178.535 ;
        RECT 109.120 178.515 109.230 178.535 ;
        RECT 107.240 178.375 107.360 178.485 ;
        RECT 108.620 178.375 108.740 178.485 ;
        RECT 109.060 178.345 109.255 178.515 ;
        RECT 109.555 178.370 109.715 178.480 ;
        RECT 113.695 178.380 113.855 178.490 ;
        RECT 109.085 178.325 109.255 178.345 ;
        RECT 114.140 178.345 114.310 178.515 ;
        RECT 114.140 178.325 114.195 178.345 ;
        RECT 115.525 178.325 115.695 178.535 ;
        RECT 41.785 177.515 43.155 178.325 ;
        RECT 43.165 177.515 48.675 178.325 ;
        RECT 49.605 177.415 52.355 178.325 ;
        RECT 52.365 177.515 57.875 178.325 ;
        RECT 58.345 177.645 62.245 178.325 ;
        RECT 62.485 177.645 65.225 178.325 ;
        RECT 58.345 177.415 59.275 177.645 ;
        RECT 65.245 177.515 67.075 178.325 ;
        RECT 68.105 177.415 70.295 178.325 ;
        RECT 70.305 177.515 75.815 178.325 ;
        RECT 75.825 177.645 79.725 178.325 ;
        RECT 79.965 178.075 85.060 178.325 ;
        RECT 87.855 178.155 89.615 178.325 ;
        RECT 87.360 178.110 89.615 178.155 ;
        RECT 86.420 178.075 89.615 178.110 ;
        RECT 79.965 177.645 89.615 178.075 ;
        RECT 75.825 177.415 76.755 177.645 ;
        RECT 79.965 177.415 81.985 177.645 ;
        RECT 81.065 177.395 81.985 177.415 ;
        RECT 85.060 177.475 88.290 177.645 ;
        RECT 89.825 177.505 91.755 178.325 ;
        RECT 91.925 177.515 93.295 178.325 ;
        RECT 93.765 177.645 97.665 178.325 ;
        RECT 85.060 177.430 87.350 177.475 ;
        RECT 85.060 177.395 86.410 177.430 ;
        RECT 89.825 177.415 90.775 177.505 ;
        RECT 93.765 177.415 94.695 177.645 ;
        RECT 98.165 177.415 102.035 178.325 ;
        RECT 102.965 177.645 106.865 178.325 ;
        RECT 107.565 177.645 109.395 178.325 ;
        RECT 102.965 177.415 103.895 177.645 ;
        RECT 107.565 177.415 108.910 177.645 ;
        RECT 110.325 177.415 114.195 178.325 ;
        RECT 114.465 177.515 115.835 178.325 ;
        RECT 41.785 173.095 43.155 173.905 ;
        RECT 43.165 173.095 48.675 173.905 ;
        RECT 48.785 173.095 51.895 174.005 ;
        RECT 51.905 173.095 54.655 173.905 ;
        RECT 55.225 173.095 58.335 174.005 ;
        RECT 58.545 173.915 59.495 174.005 ;
        RECT 58.545 173.095 60.475 173.915 ;
        RECT 60.645 173.095 62.015 173.905 ;
        RECT 65.225 173.775 66.155 174.005 ;
        RECT 62.255 173.095 66.155 173.775 ;
        RECT 66.165 173.775 67.095 174.005 ;
        RECT 73.510 173.990 74.860 174.025 ;
        RECT 72.570 173.945 74.860 173.990 ;
        RECT 71.630 173.775 74.860 173.945 ;
        RECT 77.935 174.005 78.855 174.025 ;
        RECT 77.935 173.775 79.955 174.005 ;
        RECT 84.085 173.775 85.015 174.005 ;
        RECT 66.165 173.095 70.065 173.775 ;
        RECT 70.305 173.345 79.955 173.775 ;
        RECT 70.305 173.310 73.500 173.345 ;
        RECT 70.305 173.265 72.560 173.310 ;
        RECT 70.305 173.095 72.065 173.265 ;
        RECT 74.860 173.095 79.955 173.345 ;
        RECT 81.115 173.095 85.015 173.775 ;
        RECT 85.025 173.095 86.395 173.875 ;
        RECT 86.405 173.095 88.235 173.905 ;
        RECT 91.445 173.775 92.375 174.005 ;
        RECT 95.585 173.775 96.515 174.005 ;
        RECT 88.475 173.095 92.375 173.775 ;
        RECT 92.615 173.095 96.515 173.775 ;
        RECT 97.445 173.775 98.375 174.005 ;
        RECT 101.585 173.775 102.515 174.005 ;
        RECT 106.645 173.775 107.575 174.005 ;
        RECT 97.445 173.095 101.345 173.775 ;
        RECT 101.585 173.095 105.485 173.775 ;
        RECT 106.645 173.095 110.545 173.775 ;
        RECT 111.845 173.095 114.455 174.005 ;
        RECT 114.465 173.095 115.835 173.905 ;
        RECT 41.925 172.885 42.095 173.095 ;
        RECT 43.305 172.885 43.475 173.095 ;
        RECT 48.825 172.885 48.995 173.095 ;
        RECT 52.045 172.905 52.215 173.095 ;
        RECT 54.345 172.885 54.515 173.075 ;
        RECT 55.265 172.905 55.435 173.095 ;
        RECT 60.325 173.075 60.475 173.095 ;
        RECT 56.460 172.885 56.630 173.075 ;
        RECT 60.325 172.885 60.495 173.075 ;
        RECT 60.785 172.905 60.955 173.095 ;
        RECT 62.160 172.935 62.280 173.045 ;
        RECT 62.630 172.885 62.800 173.075 ;
        RECT 65.570 172.905 65.740 173.095 ;
        RECT 66.305 172.885 66.475 173.075 ;
        RECT 66.580 172.905 66.750 173.095 ;
        RECT 68.155 172.885 68.325 173.075 ;
        RECT 69.525 172.885 69.695 173.075 ;
        RECT 70.445 172.905 70.615 173.095 ;
        RECT 75.045 172.885 75.215 173.075 ;
        RECT 80.100 172.935 80.220 173.045 ;
        RECT 80.560 172.935 80.680 173.045 ;
        RECT 81.300 172.885 81.470 173.075 ;
        RECT 84.430 172.905 84.600 173.095 ;
        RECT 86.075 173.075 86.245 173.095 ;
        RECT 85.175 172.930 85.335 173.040 ;
        RECT 86.075 172.905 86.250 173.075 ;
        RECT 86.545 172.905 86.715 173.095 ;
        RECT 86.135 172.885 86.250 172.905 ;
        RECT 91.145 172.885 91.315 173.075 ;
        RECT 91.790 172.905 91.960 173.095 ;
        RECT 92.980 172.935 93.100 173.045 ;
        RECT 93.905 172.885 94.075 173.075 ;
        RECT 95.930 172.905 96.100 173.095 ;
        RECT 96.675 173.045 96.835 173.050 ;
        RECT 96.660 172.940 96.835 173.045 ;
        RECT 96.660 172.935 96.780 172.940 ;
        RECT 97.120 172.905 97.290 173.075 ;
        RECT 97.860 172.905 98.030 173.095 ;
        RECT 102.000 172.905 102.170 173.095 ;
        RECT 97.175 172.885 97.290 172.905 ;
        RECT 102.185 172.885 102.355 173.075 ;
        RECT 104.945 172.885 105.115 173.075 ;
        RECT 105.860 172.935 105.980 173.045 ;
        RECT 107.060 172.905 107.230 173.095 ;
        RECT 110.935 172.940 111.095 173.050 ;
        RECT 114.140 172.905 114.310 173.095 ;
        RECT 115.525 172.885 115.695 173.095 ;
        RECT 41.785 172.075 43.155 172.885 ;
        RECT 43.165 172.075 48.675 172.885 ;
        RECT 48.685 172.075 54.195 172.885 ;
        RECT 54.205 172.075 56.035 172.885 ;
        RECT 56.045 172.205 59.945 172.885 ;
        RECT 56.045 171.975 56.975 172.205 ;
        RECT 60.185 172.075 62.015 172.885 ;
        RECT 62.485 172.205 66.155 172.885 ;
        RECT 65.130 171.975 66.155 172.205 ;
        RECT 66.165 172.075 67.535 172.885 ;
        RECT 68.005 172.105 69.375 172.885 ;
        RECT 69.385 172.075 74.895 172.885 ;
        RECT 74.905 172.075 80.415 172.885 ;
        RECT 80.885 172.205 84.785 172.885 ;
        RECT 80.885 171.975 81.815 172.205 ;
        RECT 86.135 171.975 90.995 172.885 ;
        RECT 91.005 172.075 92.835 172.885 ;
        RECT 93.765 172.075 96.515 172.885 ;
        RECT 97.175 171.975 102.035 172.885 ;
        RECT 102.045 172.075 104.795 172.885 ;
        RECT 104.805 172.715 106.565 172.885 ;
        RECT 104.805 172.670 107.060 172.715 ;
        RECT 104.805 172.635 108.000 172.670 ;
        RECT 109.360 172.635 114.455 172.885 ;
        RECT 104.805 172.205 114.455 172.635 ;
        RECT 106.130 172.035 109.360 172.205 ;
        RECT 107.070 171.990 109.360 172.035 ;
        RECT 108.010 171.955 109.360 171.990 ;
        RECT 112.435 171.975 114.455 172.205 ;
        RECT 114.465 172.075 115.835 172.885 ;
        RECT 112.435 171.955 113.355 171.975 ;
        RECT 41.785 167.655 43.155 168.465 ;
        RECT 43.165 167.655 48.675 168.465 ;
        RECT 48.685 167.655 54.195 168.465 ;
        RECT 55.125 167.655 58.795 168.465 ;
        RECT 58.805 167.655 60.175 168.465 ;
        RECT 63.385 168.335 64.315 168.565 ;
        RECT 60.415 167.655 64.315 168.335 ;
        RECT 64.325 167.655 67.075 168.465 ;
        RECT 70.260 168.335 71.675 168.565 ;
        RECT 67.645 167.655 71.675 168.335 ;
        RECT 71.685 168.335 72.615 168.565 ;
        RECT 85.010 168.550 86.360 168.585 ;
        RECT 84.070 168.505 86.360 168.550 ;
        RECT 71.685 167.655 75.585 168.335 ;
        RECT 75.825 167.655 79.495 168.465 ;
        RECT 83.130 168.335 86.360 168.505 ;
        RECT 89.435 168.565 90.355 168.585 ;
        RECT 89.435 168.335 91.455 168.565 ;
        RECT 95.100 168.335 96.515 168.565 ;
        RECT 99.730 168.550 101.080 168.585 ;
        RECT 98.790 168.505 101.080 168.550 ;
        RECT 97.850 168.335 101.080 168.505 ;
        RECT 104.155 168.565 105.075 168.585 ;
        RECT 104.155 168.335 106.175 168.565 ;
        RECT 81.805 167.905 91.455 168.335 ;
        RECT 81.805 167.870 85.000 167.905 ;
        RECT 81.805 167.825 84.060 167.870 ;
        RECT 81.805 167.655 83.565 167.825 ;
        RECT 86.360 167.655 91.455 167.905 ;
        RECT 92.485 167.655 96.515 168.335 ;
        RECT 96.525 167.905 106.175 168.335 ;
        RECT 96.525 167.870 99.720 167.905 ;
        RECT 96.525 167.825 98.780 167.870 ;
        RECT 96.525 167.655 98.285 167.825 ;
        RECT 101.080 167.655 106.175 167.905 ;
        RECT 106.645 168.335 107.575 168.565 ;
        RECT 106.645 167.655 110.545 168.335 ;
        RECT 110.785 167.655 112.155 168.435 ;
        RECT 112.165 167.655 113.535 168.435 ;
        RECT 114.465 167.655 115.835 168.465 ;
        RECT 41.925 167.445 42.095 167.655 ;
        RECT 43.305 167.445 43.475 167.655 ;
        RECT 48.825 167.445 48.995 167.655 ;
        RECT 54.340 167.495 54.460 167.605 ;
        RECT 55.265 167.465 55.435 167.655 ;
        RECT 58.945 167.465 59.115 167.655 ;
        RECT 59.865 167.445 60.035 167.635 ;
        RECT 60.325 167.445 60.495 167.635 ;
        RECT 63.730 167.465 63.900 167.655 ;
        RECT 64.465 167.465 64.635 167.655 ;
        RECT 65.845 167.445 66.015 167.635 ;
        RECT 67.220 167.495 67.340 167.605 ;
        RECT 67.685 167.465 67.855 167.655 ;
        RECT 68.145 167.445 68.315 167.635 ;
        RECT 72.100 167.465 72.270 167.655 ;
        RECT 72.285 167.445 72.455 167.635 ;
        RECT 72.745 167.445 72.915 167.635 ;
        RECT 74.590 167.445 74.760 167.635 ;
        RECT 75.965 167.465 76.135 167.655 ;
        RECT 78.265 167.445 78.435 167.635 ;
        RECT 79.655 167.500 79.815 167.610 ;
        RECT 81.025 167.445 81.195 167.635 ;
        RECT 81.485 167.445 81.655 167.635 ;
        RECT 81.945 167.465 82.115 167.655 ;
        RECT 87.005 167.445 87.175 167.635 ;
        RECT 90.695 167.490 90.855 167.600 ;
        RECT 91.615 167.500 91.775 167.610 ;
        RECT 92.525 167.465 92.695 167.655 ;
        RECT 92.985 167.445 93.155 167.635 ;
        RECT 93.905 167.445 94.075 167.635 ;
        RECT 96.665 167.465 96.835 167.655 ;
        RECT 98.045 167.445 98.215 167.635 ;
        RECT 103.575 167.490 103.735 167.600 ;
        RECT 107.060 167.465 107.230 167.655 ;
        RECT 109.090 167.465 109.260 167.635 ;
        RECT 109.540 167.495 109.660 167.605 ;
        RECT 109.090 167.445 109.205 167.465 ;
        RECT 110.280 167.445 110.450 167.635 ;
        RECT 111.845 167.465 112.015 167.655 ;
        RECT 113.215 167.465 113.385 167.655 ;
        RECT 113.695 167.500 113.855 167.610 ;
        RECT 114.140 167.495 114.260 167.605 ;
        RECT 115.525 167.445 115.695 167.655 ;
        RECT 41.785 166.635 43.155 167.445 ;
        RECT 43.165 166.635 48.675 167.445 ;
        RECT 48.685 166.635 50.515 167.445 ;
        RECT 50.525 167.195 55.620 167.445 ;
        RECT 58.415 167.275 60.175 167.445 ;
        RECT 57.920 167.230 60.175 167.275 ;
        RECT 56.980 167.195 60.175 167.230 ;
        RECT 50.525 166.765 60.175 167.195 ;
        RECT 50.525 166.535 52.545 166.765 ;
        RECT 51.625 166.515 52.545 166.535 ;
        RECT 55.620 166.595 58.850 166.765 ;
        RECT 60.185 166.635 65.695 167.445 ;
        RECT 65.705 166.635 67.535 167.445 ;
        RECT 68.005 166.635 70.755 167.445 ;
        RECT 70.765 166.765 72.595 167.445 ;
        RECT 72.605 166.635 74.435 167.445 ;
        RECT 74.445 166.765 78.115 167.445 ;
        RECT 55.620 166.550 57.910 166.595 ;
        RECT 55.620 166.515 56.970 166.550 ;
        RECT 77.090 166.535 78.115 166.765 ;
        RECT 78.125 166.635 79.495 167.445 ;
        RECT 79.505 166.765 81.335 167.445 ;
        RECT 81.345 166.635 86.855 167.445 ;
        RECT 86.865 166.635 90.535 167.445 ;
        RECT 91.465 166.765 93.295 167.445 ;
        RECT 93.865 166.765 97.895 167.445 ;
        RECT 96.480 166.535 97.895 166.765 ;
        RECT 97.905 166.635 103.415 167.445 ;
        RECT 104.345 166.535 109.205 167.445 ;
        RECT 109.865 166.765 113.765 167.445 ;
        RECT 109.865 166.535 110.795 166.765 ;
        RECT 114.465 166.635 115.835 167.445 ;
        RECT 62.205 163.125 63.125 163.145 ;
        RECT 41.785 162.215 43.155 163.025 ;
        RECT 43.165 162.215 48.675 163.025 ;
        RECT 48.685 162.215 54.195 163.025 ;
        RECT 55.125 162.215 58.235 163.125 ;
        RECT 58.345 162.215 61.095 163.025 ;
        RECT 61.105 162.895 63.125 163.125 ;
        RECT 66.200 163.110 67.550 163.145 ;
        RECT 66.200 163.065 68.490 163.110 ;
        RECT 66.200 162.895 69.430 163.065 ;
        RECT 61.105 162.465 70.755 162.895 ;
        RECT 61.105 162.215 66.200 162.465 ;
        RECT 67.560 162.430 70.755 162.465 ;
        RECT 68.500 162.385 70.755 162.430 ;
        RECT 68.995 162.215 70.755 162.385 ;
        RECT 70.765 162.215 76.275 163.025 ;
        RECT 76.285 162.215 78.115 163.025 ;
        RECT 83.600 162.895 85.015 163.125 ;
        RECT 78.585 162.215 80.415 162.895 ;
        RECT 80.985 162.215 85.015 162.895 ;
        RECT 85.945 162.895 86.875 163.125 ;
        RECT 85.945 162.215 89.845 162.895 ;
        RECT 90.085 162.215 93.755 163.025 ;
        RECT 93.765 162.895 94.695 163.125 ;
        RECT 97.905 162.895 98.835 163.125 ;
        RECT 93.765 162.215 97.665 162.895 ;
        RECT 97.905 162.215 101.805 162.895 ;
        RECT 102.045 162.215 103.875 162.895 ;
        RECT 103.885 162.215 105.715 163.025 ;
        RECT 106.645 162.215 109.395 163.025 ;
        RECT 109.405 162.215 110.775 162.995 ;
        RECT 110.785 162.215 112.155 162.995 ;
        RECT 112.165 162.215 113.535 162.995 ;
        RECT 114.465 162.215 115.835 163.025 ;
        RECT 41.925 162.005 42.095 162.215 ;
        RECT 43.305 162.005 43.475 162.215 ;
        RECT 48.825 162.005 48.995 162.215 ;
        RECT 51.580 162.055 51.700 162.165 ;
        RECT 52.045 162.005 52.215 162.195 ;
        RECT 54.340 162.055 54.460 162.165 ;
        RECT 55.265 162.005 55.435 162.195 ;
        RECT 58.025 162.025 58.195 162.215 ;
        RECT 58.485 162.005 58.655 162.215 ;
        RECT 61.245 162.005 61.415 162.195 ;
        RECT 64.465 162.005 64.635 162.195 ;
        RECT 68.145 162.005 68.315 162.195 ;
        RECT 70.260 162.005 70.430 162.195 ;
        RECT 70.445 162.025 70.615 162.215 ;
        RECT 70.905 162.025 71.075 162.215 ;
        RECT 74.400 162.005 74.570 162.195 ;
        RECT 76.425 162.025 76.595 162.215 ;
        RECT 78.260 162.160 78.380 162.165 ;
        RECT 78.260 162.055 78.435 162.160 ;
        RECT 78.275 162.050 78.435 162.055 ;
        RECT 79.185 162.005 79.355 162.195 ;
        RECT 80.105 162.025 80.275 162.215 ;
        RECT 81.025 162.025 81.195 162.215 ;
        RECT 82.405 162.005 82.575 162.195 ;
        RECT 85.175 162.060 85.335 162.170 ;
        RECT 86.360 162.025 86.530 162.215 ;
        RECT 87.925 162.005 88.095 162.195 ;
        RECT 90.225 162.025 90.395 162.215 ;
        RECT 92.525 162.005 92.695 162.195 ;
        RECT 92.980 162.055 93.100 162.165 ;
        RECT 93.905 162.005 94.075 162.195 ;
        RECT 94.180 162.025 94.350 162.215 ;
        RECT 97.125 162.005 97.295 162.195 ;
        RECT 97.585 162.005 97.755 162.195 ;
        RECT 98.320 162.025 98.490 162.215 ;
        RECT 101.260 162.055 101.380 162.165 ;
        RECT 102.000 162.005 102.170 162.195 ;
        RECT 102.185 162.025 102.355 162.215 ;
        RECT 104.025 162.025 104.195 162.215 ;
        RECT 105.860 162.055 105.980 162.165 ;
        RECT 106.785 162.025 106.955 162.215 ;
        RECT 109.080 162.005 109.250 162.195 ;
        RECT 109.545 162.005 109.715 162.195 ;
        RECT 110.455 162.025 110.625 162.215 ;
        RECT 111.845 162.195 112.015 162.215 ;
        RECT 111.835 162.025 112.015 162.195 ;
        RECT 111.835 162.005 112.005 162.025 ;
        RECT 113.225 162.005 113.395 162.215 ;
        RECT 113.695 162.050 113.855 162.170 ;
        RECT 115.525 162.005 115.695 162.215 ;
        RECT 41.785 161.195 43.155 162.005 ;
        RECT 43.165 161.195 48.675 162.005 ;
        RECT 48.685 161.195 51.435 162.005 ;
        RECT 51.945 161.095 55.115 162.005 ;
        RECT 55.225 161.095 58.335 162.005 ;
        RECT 58.345 161.195 61.095 162.005 ;
        RECT 61.205 161.095 64.315 162.005 ;
        RECT 64.365 161.095 67.535 162.005 ;
        RECT 68.005 161.195 69.835 162.005 ;
        RECT 69.845 161.325 73.745 162.005 ;
        RECT 73.985 161.325 77.885 162.005 ;
        RECT 69.845 161.095 70.775 161.325 ;
        RECT 73.985 161.095 74.915 161.325 ;
        RECT 79.145 161.095 82.255 162.005 ;
        RECT 82.265 161.195 87.775 162.005 ;
        RECT 87.785 161.195 89.615 162.005 ;
        RECT 89.625 161.095 92.795 162.005 ;
        RECT 93.765 161.195 95.595 162.005 ;
        RECT 95.605 161.325 97.435 162.005 ;
        RECT 97.445 161.195 101.115 162.005 ;
        RECT 101.585 161.325 105.485 162.005 ;
        RECT 105.725 161.325 109.395 162.005 ;
        RECT 101.585 161.095 102.515 161.325 ;
        RECT 105.725 161.095 106.750 161.325 ;
        RECT 109.405 161.195 110.775 162.005 ;
        RECT 110.785 161.225 112.155 162.005 ;
        RECT 112.165 161.225 113.535 162.005 ;
        RECT 114.465 161.195 115.835 162.005 ;
        RECT 41.785 156.775 43.155 157.585 ;
        RECT 43.625 156.775 44.995 157.555 ;
        RECT 45.005 156.775 48.675 157.585 ;
        RECT 48.685 156.775 50.055 157.555 ;
        RECT 50.065 156.775 53.735 157.585 ;
        RECT 55.125 156.775 56.495 157.555 ;
        RECT 56.505 156.775 58.335 157.585 ;
        RECT 58.805 156.775 60.175 157.555 ;
        RECT 60.185 156.775 63.855 157.585 ;
        RECT 63.865 156.775 65.235 157.555 ;
        RECT 65.245 156.775 67.075 157.585 ;
        RECT 68.105 156.775 71.215 157.685 ;
        RECT 71.225 156.775 72.595 157.555 ;
        RECT 72.605 156.775 73.975 157.585 ;
        RECT 73.985 156.775 75.355 157.555 ;
        RECT 75.365 156.775 79.035 157.585 ;
        RECT 79.045 156.775 80.415 157.555 ;
        RECT 80.885 156.775 82.715 157.585 ;
        RECT 83.185 156.775 86.295 157.685 ;
        RECT 86.405 156.775 87.775 157.555 ;
        RECT 87.785 156.775 89.155 157.585 ;
        RECT 89.165 156.775 90.535 157.555 ;
        RECT 90.545 156.775 93.295 157.585 ;
        RECT 94.225 156.775 95.595 157.555 ;
        RECT 95.605 156.775 99.275 157.585 ;
        RECT 99.285 156.775 100.655 157.555 ;
        RECT 100.665 156.775 104.335 157.585 ;
        RECT 104.345 156.775 105.715 157.555 ;
        RECT 109.360 157.455 110.775 157.685 ;
        RECT 106.745 156.775 110.775 157.455 ;
        RECT 110.785 156.775 112.155 157.555 ;
        RECT 113.085 156.775 114.455 157.555 ;
        RECT 114.465 156.775 115.835 157.585 ;
        RECT 41.925 156.585 42.095 156.775 ;
        RECT 43.300 156.615 43.420 156.725 ;
        RECT 43.775 156.585 43.945 156.775 ;
        RECT 45.145 156.585 45.315 156.775 ;
        RECT 48.835 156.585 49.005 156.775 ;
        RECT 50.205 156.585 50.375 156.775 ;
        RECT 53.895 156.620 54.055 156.730 ;
        RECT 55.275 156.585 55.445 156.775 ;
        RECT 56.645 156.585 56.815 156.775 ;
        RECT 58.480 156.615 58.600 156.725 ;
        RECT 58.945 156.585 59.115 156.775 ;
        RECT 60.325 156.585 60.495 156.775 ;
        RECT 64.015 156.585 64.185 156.775 ;
        RECT 65.385 156.585 65.555 156.775 ;
        RECT 67.220 156.615 67.340 156.725 ;
        RECT 68.145 156.585 68.315 156.775 ;
        RECT 71.365 156.585 71.535 156.775 ;
        RECT 72.745 156.585 72.915 156.775 ;
        RECT 74.135 156.585 74.305 156.775 ;
        RECT 75.505 156.585 75.675 156.775 ;
        RECT 80.095 156.585 80.265 156.775 ;
        RECT 81.025 156.585 81.195 156.775 ;
        RECT 82.860 156.615 82.980 156.725 ;
        RECT 86.085 156.585 86.255 156.775 ;
        RECT 86.555 156.585 86.725 156.775 ;
        RECT 87.925 156.585 88.095 156.775 ;
        RECT 89.305 156.585 89.475 156.775 ;
        RECT 90.685 156.585 90.855 156.775 ;
        RECT 93.900 156.615 94.020 156.725 ;
        RECT 94.375 156.585 94.545 156.775 ;
        RECT 95.745 156.585 95.915 156.775 ;
        RECT 99.425 156.585 99.595 156.775 ;
        RECT 100.805 156.585 100.975 156.775 ;
        RECT 104.495 156.585 104.665 156.775 ;
        RECT 105.860 156.615 105.980 156.725 ;
        RECT 106.785 156.585 106.955 156.775 ;
        RECT 110.935 156.585 111.105 156.775 ;
        RECT 112.315 156.620 112.475 156.730 ;
        RECT 114.135 156.585 114.305 156.775 ;
        RECT 115.525 156.585 115.695 156.775 ;
        RECT 78.050 111.500 80.060 127.610 ;
        RECT 100.710 111.500 102.720 127.610 ;
        RECT 123.370 111.500 125.380 127.610 ;
        RECT 55.390 94.160 57.400 110.270 ;
        RECT 78.050 94.160 80.060 110.270 ;
        RECT 100.710 94.160 102.720 110.270 ;
        RECT 123.370 94.160 125.380 110.270 ;
        RECT 55.390 76.820 57.400 92.930 ;
        RECT 78.050 76.820 80.060 92.930 ;
        RECT 100.710 76.820 102.720 92.930 ;
        RECT 123.370 76.820 125.380 92.930 ;
        RECT 55.390 59.480 57.400 75.590 ;
        RECT 78.050 59.480 80.060 75.590 ;
        RECT 100.710 59.480 102.720 75.590 ;
        RECT 123.370 59.480 125.380 75.590 ;
      LAYER li1 ;
        RECT 44.165 185.535 44.475 186.335 ;
        RECT 47.935 185.575 48.105 186.335 ;
        RECT 50.235 185.575 50.405 186.335 ;
        RECT 52.075 185.575 52.245 186.335 ;
        RECT 56.615 185.575 56.785 186.335 ;
        RECT 44.165 185.365 45.195 185.535 ;
        RECT 47.935 185.405 48.650 185.575 ;
        RECT 50.235 185.405 50.950 185.575 ;
        RECT 52.075 185.405 52.790 185.575 ;
        RECT 44.165 184.455 44.335 185.365 ;
        RECT 45.025 185.115 45.195 185.365 ;
        RECT 48.480 185.195 48.650 185.405 ;
        RECT 50.780 185.195 50.950 185.405 ;
        RECT 52.620 185.195 52.790 185.405 ;
        RECT 56.070 185.405 56.785 185.575 ;
        RECT 57.595 185.575 57.765 186.335 ;
        RECT 59.435 185.575 59.605 186.335 ;
        RECT 62.595 185.575 62.765 186.335 ;
        RECT 57.595 185.405 58.310 185.575 ;
        RECT 59.435 185.405 60.150 185.575 ;
        RECT 56.070 185.195 56.240 185.405 ;
        RECT 45.025 184.945 46.165 185.115 ;
        RECT 48.480 184.865 48.735 185.195 ;
        RECT 50.780 184.865 51.035 185.195 ;
        RECT 52.620 184.865 52.875 185.195 ;
        RECT 55.985 184.865 56.240 185.195 ;
        RECT 48.480 184.675 48.650 184.865 ;
        RECT 50.780 184.675 50.950 184.865 ;
        RECT 52.620 184.675 52.790 184.865 ;
        RECT 47.935 184.505 48.650 184.675 ;
        RECT 50.235 184.505 50.950 184.675 ;
        RECT 52.075 184.505 52.790 184.675 ;
        RECT 56.070 184.675 56.240 184.865 ;
        RECT 57.505 184.855 57.860 185.225 ;
        RECT 58.140 185.195 58.310 185.405 ;
        RECT 58.140 184.865 58.395 185.195 ;
        RECT 58.140 184.675 58.310 184.865 ;
        RECT 59.345 184.855 59.700 185.225 ;
        RECT 59.980 185.195 60.150 185.405 ;
        RECT 62.050 185.405 62.765 185.575 ;
        RECT 63.025 185.535 63.335 186.335 ;
        RECT 65.875 185.575 66.045 186.335 ;
        RECT 69.495 185.575 69.665 186.335 ;
        RECT 62.050 185.195 62.220 185.405 ;
        RECT 63.025 185.365 64.055 185.535 ;
        RECT 65.875 185.405 66.590 185.575 ;
        RECT 59.980 184.865 60.235 185.195 ;
        RECT 61.965 184.865 62.220 185.195 ;
        RECT 59.980 184.675 60.150 184.865 ;
        RECT 56.070 184.505 56.785 184.675 ;
        RECT 44.165 184.125 44.465 184.455 ;
        RECT 47.935 184.125 48.105 184.505 ;
        RECT 50.235 184.125 50.405 184.505 ;
        RECT 52.075 184.125 52.245 184.505 ;
        RECT 56.615 184.125 56.785 184.505 ;
        RECT 57.595 184.505 58.310 184.675 ;
        RECT 59.435 184.505 60.150 184.675 ;
        RECT 62.050 184.675 62.220 184.865 ;
        RECT 62.500 184.855 62.855 185.225 ;
        RECT 62.050 184.505 62.765 184.675 ;
        RECT 57.595 184.125 57.765 184.505 ;
        RECT 59.435 184.125 59.605 184.505 ;
        RECT 62.595 184.125 62.765 184.505 ;
        RECT 63.025 184.455 63.195 185.365 ;
        RECT 63.365 184.625 63.715 185.195 ;
        RECT 63.885 185.115 64.055 185.365 ;
        RECT 63.885 184.945 65.025 185.115 ;
        RECT 65.785 184.855 66.140 185.225 ;
        RECT 66.420 185.195 66.590 185.405 ;
        RECT 68.950 185.405 69.665 185.575 ;
        RECT 70.015 185.575 70.185 186.335 ;
        RECT 73.175 185.575 73.345 186.335 ;
        RECT 75.935 185.575 76.105 186.335 ;
        RECT 78.235 185.575 78.405 186.335 ;
        RECT 70.015 185.405 70.730 185.575 ;
        RECT 68.950 185.195 69.120 185.405 ;
        RECT 66.420 184.865 66.675 185.195 ;
        RECT 68.865 184.865 69.120 185.195 ;
        RECT 66.420 184.675 66.590 184.865 ;
        RECT 65.875 184.505 66.590 184.675 ;
        RECT 68.950 184.675 69.120 184.865 ;
        RECT 69.400 184.855 69.755 185.225 ;
        RECT 69.925 184.855 70.280 185.225 ;
        RECT 70.560 185.195 70.730 185.405 ;
        RECT 72.630 185.405 73.345 185.575 ;
        RECT 75.390 185.405 76.105 185.575 ;
        RECT 77.690 185.405 78.405 185.575 ;
        RECT 84.135 185.525 84.465 186.335 ;
        RECT 86.925 185.535 87.235 186.335 ;
        RECT 72.630 185.195 72.800 185.405 ;
        RECT 70.560 184.865 70.815 185.195 ;
        RECT 72.545 184.865 72.800 185.195 ;
        RECT 70.560 184.675 70.730 184.865 ;
        RECT 68.950 184.505 69.665 184.675 ;
        RECT 63.025 184.125 63.325 184.455 ;
        RECT 65.875 184.125 66.045 184.505 ;
        RECT 69.495 184.125 69.665 184.505 ;
        RECT 70.015 184.505 70.730 184.675 ;
        RECT 72.630 184.675 72.800 184.865 ;
        RECT 73.080 184.855 73.435 185.225 ;
        RECT 75.390 185.195 75.560 185.405 ;
        RECT 75.305 184.865 75.560 185.195 ;
        RECT 75.390 184.675 75.560 184.865 ;
        RECT 75.840 184.855 76.195 185.225 ;
        RECT 77.690 185.195 77.860 185.405 ;
        RECT 83.750 185.355 84.465 185.525 ;
        RECT 86.205 185.365 87.235 185.535 ;
        RECT 77.605 184.865 77.860 185.195 ;
        RECT 77.690 184.675 77.860 184.865 ;
        RECT 78.140 184.855 78.495 185.225 ;
        RECT 83.750 185.115 83.920 185.355 ;
        RECT 83.420 184.945 83.920 185.115 ;
        RECT 84.090 184.945 84.470 185.185 ;
        RECT 86.205 185.115 86.375 185.365 ;
        RECT 85.235 184.945 86.375 185.115 ;
        RECT 83.750 184.775 83.920 184.945 ;
        RECT 72.630 184.505 73.345 184.675 ;
        RECT 75.390 184.505 76.105 184.675 ;
        RECT 77.690 184.505 78.405 184.675 ;
        RECT 83.750 184.605 84.385 184.775 ;
        RECT 86.545 184.625 86.895 185.195 ;
        RECT 70.015 184.125 70.185 184.505 ;
        RECT 73.175 184.125 73.345 184.505 ;
        RECT 75.935 184.125 76.105 184.505 ;
        RECT 78.235 184.125 78.405 184.505 ;
        RECT 84.215 184.125 84.385 184.605 ;
        RECT 87.065 184.455 87.235 185.365 ;
        RECT 86.935 184.125 87.235 184.455 ;
        RECT 87.405 185.430 87.675 186.335 ;
        RECT 88.355 185.575 88.535 186.335 ;
        RECT 87.405 184.630 87.585 185.430 ;
        RECT 87.860 185.405 88.535 185.575 ;
        RECT 89.245 185.430 89.515 186.335 ;
        RECT 90.195 185.575 90.365 186.335 ;
        RECT 87.860 185.260 88.030 185.405 ;
        RECT 87.755 184.930 88.030 185.260 ;
        RECT 87.860 184.675 88.030 184.930 ;
        RECT 87.405 184.125 87.665 184.630 ;
        RECT 87.860 184.505 88.525 184.675 ;
        RECT 88.355 184.125 88.525 184.505 ;
        RECT 89.245 184.630 89.415 185.430 ;
        RECT 89.700 185.405 90.365 185.575 ;
        RECT 91.085 185.430 91.355 186.335 ;
        RECT 92.035 185.575 92.215 186.335 ;
        RECT 89.700 185.260 89.870 185.405 ;
        RECT 89.585 184.930 89.870 185.260 ;
        RECT 89.700 184.675 89.870 184.930 ;
        RECT 89.245 184.125 89.505 184.630 ;
        RECT 89.700 184.505 90.365 184.675 ;
        RECT 90.195 184.125 90.365 184.505 ;
        RECT 91.085 184.630 91.265 185.430 ;
        RECT 91.540 185.405 92.215 185.575 ;
        RECT 96.795 185.525 97.125 186.335 ;
        RECT 101.185 185.535 101.495 186.335 ;
        RECT 102.755 186.165 104.785 186.335 ;
        RECT 91.540 185.260 91.710 185.405 ;
        RECT 91.435 184.930 91.710 185.260 ;
        RECT 96.375 185.355 97.125 185.525 ;
        RECT 100.465 185.365 101.495 185.535 ;
        RECT 96.375 185.115 96.545 185.355 ;
        RECT 96.075 184.945 96.545 185.115 ;
        RECT 96.715 184.945 97.620 185.185 ;
        RECT 100.465 185.115 100.635 185.365 ;
        RECT 99.495 184.945 100.635 185.115 ;
        RECT 91.540 184.675 91.710 184.930 ;
        RECT 96.375 184.775 96.545 184.945 ;
        RECT 91.085 184.125 91.345 184.630 ;
        RECT 91.540 184.505 92.205 184.675 ;
        RECT 96.375 184.605 97.125 184.775 ;
        RECT 100.805 184.625 101.155 185.195 ;
        RECT 92.035 184.125 92.205 184.505 ;
        RECT 96.795 184.125 97.125 184.605 ;
        RECT 101.325 184.455 101.495 185.365 ;
        RECT 101.665 185.745 102.180 186.155 ;
        RECT 101.665 184.935 102.005 185.745 ;
        RECT 102.755 185.500 102.925 186.165 ;
        RECT 103.320 185.825 104.445 185.995 ;
        RECT 102.175 185.310 102.925 185.500 ;
        RECT 103.095 185.485 104.105 185.655 ;
        RECT 101.665 184.765 102.895 184.935 ;
        RECT 101.195 184.125 101.495 184.455 ;
        RECT 101.940 184.160 102.185 184.765 ;
        RECT 103.095 184.125 103.285 185.485 ;
        RECT 103.455 184.465 103.730 185.285 ;
        RECT 103.935 184.685 104.105 185.485 ;
        RECT 104.275 184.695 104.445 185.825 ;
        RECT 104.615 185.195 104.785 186.165 ;
        RECT 105.295 185.365 105.630 186.335 ;
        RECT 104.615 184.865 104.810 185.195 ;
        RECT 105.035 184.865 105.290 185.195 ;
        RECT 105.035 184.695 105.205 184.865 ;
        RECT 105.460 184.695 105.630 185.365 ;
        RECT 104.275 184.525 105.205 184.695 ;
        RECT 104.275 184.490 104.450 184.525 ;
        RECT 103.455 184.295 103.735 184.465 ;
        RECT 103.455 184.125 103.730 184.295 ;
        RECT 103.920 184.125 104.450 184.490 ;
        RECT 105.375 184.125 105.630 184.695 ;
        RECT 108.085 185.430 108.340 186.335 ;
        RECT 109.055 185.575 109.225 186.335 ;
        RECT 108.085 184.700 108.255 185.430 ;
        RECT 108.510 185.405 109.225 185.575 ;
        RECT 108.510 185.195 108.680 185.405 ;
        RECT 108.425 184.865 108.680 185.195 ;
        RECT 108.085 184.125 108.340 184.700 ;
        RECT 108.510 184.675 108.680 184.865 ;
        RECT 109.490 185.365 109.825 186.335 ;
        RECT 110.335 186.165 112.365 186.335 ;
        RECT 109.490 184.695 109.660 185.365 ;
        RECT 110.335 185.195 110.505 186.165 ;
        RECT 109.830 184.865 110.085 185.195 ;
        RECT 110.310 184.865 110.505 185.195 ;
        RECT 110.675 185.825 111.800 185.995 ;
        RECT 109.915 184.695 110.085 184.865 ;
        RECT 110.675 184.695 110.845 185.825 ;
        RECT 108.510 184.505 109.225 184.675 ;
        RECT 109.055 184.125 109.225 184.505 ;
        RECT 109.490 184.125 109.745 184.695 ;
        RECT 109.915 184.525 110.845 184.695 ;
        RECT 111.015 185.485 112.025 185.655 ;
        RECT 111.015 184.685 111.185 185.485 ;
        RECT 110.670 184.490 110.845 184.525 ;
        RECT 110.670 184.125 111.200 184.490 ;
        RECT 111.390 184.465 111.665 185.285 ;
        RECT 111.385 184.295 111.665 184.465 ;
        RECT 111.390 184.125 111.665 184.295 ;
        RECT 111.835 184.125 112.025 185.485 ;
        RECT 112.195 185.500 112.365 186.165 ;
        RECT 112.940 185.745 113.455 186.155 ;
        RECT 112.195 185.310 112.945 185.500 ;
        RECT 113.115 184.935 113.455 185.745 ;
        RECT 112.225 184.765 113.455 184.935 ;
        RECT 112.935 184.160 113.180 184.765 ;
        RECT 45.575 183.235 45.745 183.615 ;
        RECT 45.030 183.065 45.745 183.235 ;
        RECT 46.095 183.235 46.265 183.615 ;
        RECT 46.095 183.065 46.810 183.235 ;
        RECT 45.030 182.875 45.200 183.065 ;
        RECT 44.945 182.545 45.200 182.875 ;
        RECT 45.030 182.335 45.200 182.545 ;
        RECT 46.640 182.875 46.810 183.065 ;
        RECT 53.795 182.965 54.125 183.385 ;
        RECT 54.305 183.300 55.095 183.565 ;
        RECT 53.875 182.875 54.125 182.965 ;
        RECT 46.640 182.545 46.895 182.875 ;
        RECT 46.640 182.335 46.810 182.545 ;
        RECT 45.030 182.165 45.745 182.335 ;
        RECT 45.575 181.405 45.745 182.165 ;
        RECT 46.095 182.165 46.810 182.335 ;
        RECT 46.095 181.405 46.265 182.165 ;
        RECT 53.365 181.915 53.705 182.795 ;
        RECT 53.875 182.625 54.670 182.875 ;
        RECT 53.875 181.405 54.045 182.625 ;
        RECT 54.840 182.445 55.095 183.300 ;
        RECT 55.265 183.145 55.465 183.565 ;
        RECT 55.265 182.625 55.675 183.145 ;
        RECT 56.155 183.135 56.415 183.615 ;
        RECT 55.845 182.445 56.075 182.875 ;
        RECT 54.285 182.275 56.075 182.445 ;
        RECT 54.285 181.910 54.535 182.275 ;
        RECT 55.255 181.980 55.970 182.275 ;
        RECT 56.245 182.105 56.415 183.135 ;
        RECT 56.600 183.235 56.875 183.375 ;
        RECT 57.545 183.235 57.755 183.405 ;
        RECT 56.600 183.045 57.755 183.235 ;
        RECT 57.925 183.235 58.255 183.615 ;
        RECT 57.925 183.030 58.775 183.235 ;
        RECT 56.595 182.420 56.855 182.875 ;
        RECT 57.110 182.470 57.695 182.845 ;
        RECT 55.070 181.405 55.545 181.745 ;
        RECT 56.140 181.405 56.415 182.105 ;
        RECT 57.110 182.085 57.315 182.470 ;
        RECT 57.865 182.255 58.275 182.860 ;
        RECT 58.445 182.540 58.775 183.030 ;
        RECT 63.760 182.975 64.005 183.580 ;
        RECT 63.485 182.805 64.715 182.975 ;
        RECT 58.445 182.085 58.615 182.540 ;
        RECT 57.105 181.915 57.315 182.085 ;
        RECT 57.110 181.885 57.315 181.915 ;
        RECT 57.495 181.865 58.615 182.085 ;
        RECT 63.485 181.995 63.825 182.805 ;
        RECT 63.995 182.240 64.745 182.430 ;
        RECT 57.495 181.405 57.755 181.865 ;
        RECT 63.485 181.585 64.000 181.995 ;
        RECT 64.575 181.575 64.745 182.240 ;
        RECT 64.915 182.255 65.105 183.615 ;
        RECT 65.275 182.765 65.550 183.615 ;
        RECT 65.740 183.250 66.270 183.615 ;
        RECT 66.095 183.215 66.270 183.250 ;
        RECT 65.275 182.595 65.555 182.765 ;
        RECT 65.275 182.455 65.550 182.595 ;
        RECT 65.755 182.255 65.925 183.055 ;
        RECT 64.915 182.085 65.925 182.255 ;
        RECT 66.095 183.045 67.025 183.215 ;
        RECT 67.195 183.045 67.450 183.615 ;
        RECT 66.095 181.915 66.265 183.045 ;
        RECT 66.855 182.875 67.025 183.045 ;
        RECT 65.140 181.745 66.265 181.915 ;
        RECT 66.435 182.545 66.630 182.875 ;
        RECT 66.855 182.545 67.110 182.875 ;
        RECT 66.435 181.575 66.605 182.545 ;
        RECT 67.280 182.375 67.450 183.045 ;
        RECT 69.280 182.975 69.525 183.580 ;
        RECT 64.575 181.405 66.605 181.575 ;
        RECT 67.115 181.405 67.450 182.375 ;
        RECT 69.005 182.805 70.235 182.975 ;
        RECT 69.005 181.995 69.345 182.805 ;
        RECT 69.515 182.240 70.265 182.430 ;
        RECT 69.005 181.585 69.520 181.995 ;
        RECT 70.095 181.575 70.265 182.240 ;
        RECT 70.435 182.255 70.625 183.615 ;
        RECT 70.795 182.765 71.070 183.615 ;
        RECT 71.260 183.250 71.790 183.615 ;
        RECT 71.615 183.215 71.790 183.250 ;
        RECT 70.795 182.595 71.075 182.765 ;
        RECT 70.795 182.455 71.070 182.595 ;
        RECT 71.275 182.255 71.445 183.055 ;
        RECT 70.435 182.085 71.445 182.255 ;
        RECT 71.615 183.045 72.545 183.215 ;
        RECT 72.715 183.045 72.970 183.615 ;
        RECT 71.615 181.915 71.785 183.045 ;
        RECT 72.375 182.875 72.545 183.045 ;
        RECT 70.660 181.745 71.785 181.915 ;
        RECT 71.955 182.545 72.150 182.875 ;
        RECT 72.375 182.545 72.630 182.875 ;
        RECT 71.955 181.575 72.125 182.545 ;
        RECT 72.800 182.375 72.970 183.045 ;
        RECT 73.420 182.975 73.665 183.580 ;
        RECT 70.095 181.405 72.125 181.575 ;
        RECT 72.635 181.405 72.970 182.375 ;
        RECT 73.145 182.805 74.375 182.975 ;
        RECT 73.145 181.995 73.485 182.805 ;
        RECT 73.655 182.240 74.405 182.430 ;
        RECT 73.145 181.585 73.660 181.995 ;
        RECT 74.235 181.575 74.405 182.240 ;
        RECT 74.575 182.255 74.765 183.615 ;
        RECT 74.935 182.765 75.210 183.615 ;
        RECT 75.400 183.250 75.930 183.615 ;
        RECT 75.755 183.215 75.930 183.250 ;
        RECT 74.935 182.595 75.215 182.765 ;
        RECT 74.935 182.455 75.210 182.595 ;
        RECT 75.415 182.255 75.585 183.055 ;
        RECT 74.575 182.085 75.585 182.255 ;
        RECT 75.755 183.045 76.685 183.215 ;
        RECT 76.855 183.045 77.110 183.615 ;
        RECT 75.755 181.915 75.925 183.045 ;
        RECT 76.515 182.875 76.685 183.045 ;
        RECT 74.800 181.745 75.925 181.915 ;
        RECT 76.095 182.545 76.290 182.875 ;
        RECT 76.515 182.545 76.770 182.875 ;
        RECT 76.095 181.575 76.265 182.545 ;
        RECT 76.940 182.375 77.110 183.045 ;
        RECT 74.235 181.405 76.265 181.575 ;
        RECT 76.775 181.405 77.110 182.375 ;
        RECT 77.285 183.045 77.545 183.615 ;
        RECT 78.270 183.215 78.525 183.615 ;
        RECT 77.715 183.045 78.525 183.215 ;
        RECT 78.715 183.045 78.960 183.615 ;
        RECT 79.685 183.215 79.940 183.615 ;
        RECT 79.130 183.045 79.940 183.215 ;
        RECT 80.130 183.045 80.555 183.615 ;
        RECT 81.280 183.215 81.715 183.615 ;
        RECT 80.725 183.045 81.715 183.215 ;
        RECT 81.890 183.045 82.145 183.615 ;
        RECT 83.070 183.250 83.600 183.615 ;
        RECT 83.070 183.215 83.245 183.250 ;
        RECT 82.315 183.045 83.245 183.215 ;
        RECT 77.285 182.375 77.470 183.045 ;
        RECT 77.715 182.875 78.065 183.045 ;
        RECT 78.715 182.875 78.885 183.045 ;
        RECT 79.130 182.875 79.480 183.045 ;
        RECT 80.130 182.875 80.480 183.045 ;
        RECT 80.725 182.875 81.060 183.045 ;
        RECT 77.640 182.545 78.065 182.875 ;
        RECT 77.285 181.405 77.545 182.375 ;
        RECT 77.715 182.025 78.065 182.545 ;
        RECT 78.235 182.375 78.885 182.875 ;
        RECT 79.055 182.545 79.480 182.875 ;
        RECT 78.235 182.195 78.960 182.375 ;
        RECT 77.715 181.830 78.525 182.025 ;
        RECT 78.270 181.405 78.525 181.830 ;
        RECT 78.715 181.405 78.960 182.195 ;
        RECT 79.130 182.025 79.480 182.545 ;
        RECT 79.650 182.375 80.480 182.875 ;
        RECT 80.650 182.545 81.060 182.875 ;
        RECT 79.650 182.195 80.555 182.375 ;
        RECT 79.130 181.830 79.960 182.025 ;
        RECT 79.685 181.405 79.960 181.830 ;
        RECT 80.130 181.405 80.555 182.195 ;
        RECT 80.725 182.000 81.060 182.545 ;
        RECT 81.230 182.170 81.715 182.875 ;
        RECT 81.890 182.375 82.060 183.045 ;
        RECT 82.315 182.875 82.485 183.045 ;
        RECT 82.230 182.545 82.485 182.875 ;
        RECT 82.710 182.545 82.905 182.875 ;
        RECT 80.725 181.830 81.715 182.000 ;
        RECT 81.280 181.405 81.715 181.830 ;
        RECT 81.890 181.405 82.225 182.375 ;
        RECT 82.735 181.575 82.905 182.545 ;
        RECT 83.075 181.915 83.245 183.045 ;
        RECT 83.415 182.255 83.585 183.055 ;
        RECT 83.790 182.765 84.065 183.615 ;
        RECT 83.785 182.595 84.065 182.765 ;
        RECT 83.790 182.455 84.065 182.595 ;
        RECT 84.235 182.255 84.425 183.615 ;
        RECT 85.335 182.975 85.580 183.580 ;
        RECT 87.870 183.045 88.125 183.615 ;
        RECT 89.050 183.250 89.580 183.615 ;
        RECT 89.050 183.215 89.225 183.250 ;
        RECT 88.295 183.045 89.225 183.215 ;
        RECT 89.770 183.105 90.045 183.615 ;
        RECT 84.625 182.805 85.855 182.975 ;
        RECT 83.415 182.085 84.425 182.255 ;
        RECT 84.595 182.240 85.345 182.430 ;
        RECT 83.075 181.745 84.200 181.915 ;
        RECT 84.595 181.575 84.765 182.240 ;
        RECT 85.515 181.995 85.855 182.805 ;
        RECT 85.340 181.585 85.855 181.995 ;
        RECT 87.870 182.375 88.040 183.045 ;
        RECT 88.295 182.875 88.465 183.045 ;
        RECT 88.210 182.545 88.465 182.875 ;
        RECT 88.690 182.545 88.885 182.875 ;
        RECT 82.735 181.405 84.765 181.575 ;
        RECT 87.870 181.405 88.205 182.375 ;
        RECT 88.715 181.575 88.885 182.545 ;
        RECT 89.055 181.915 89.225 183.045 ;
        RECT 89.395 182.255 89.565 183.055 ;
        RECT 89.765 182.935 90.045 183.105 ;
        RECT 89.770 182.455 90.045 182.935 ;
        RECT 90.215 182.255 90.405 183.615 ;
        RECT 91.315 182.975 91.560 183.580 ;
        RECT 92.005 183.110 92.265 183.615 ;
        RECT 92.955 183.235 93.125 183.615 ;
        RECT 90.605 182.805 91.835 182.975 ;
        RECT 89.395 182.085 90.405 182.255 ;
        RECT 90.575 182.240 91.325 182.430 ;
        RECT 89.055 181.745 90.180 181.915 ;
        RECT 90.575 181.575 90.745 182.240 ;
        RECT 91.495 181.995 91.835 182.805 ;
        RECT 91.320 181.585 91.835 181.995 ;
        RECT 92.005 182.310 92.175 183.110 ;
        RECT 92.460 183.065 93.125 183.235 ;
        RECT 92.460 182.810 92.630 183.065 ;
        RECT 92.345 182.480 92.630 182.810 ;
        RECT 92.460 182.335 92.630 182.480 ;
        RECT 93.850 183.045 94.105 183.615 ;
        RECT 95.030 183.250 95.560 183.615 ;
        RECT 95.030 183.215 95.205 183.250 ;
        RECT 94.275 183.045 95.205 183.215 ;
        RECT 93.850 182.375 94.020 183.045 ;
        RECT 94.275 182.875 94.445 183.045 ;
        RECT 94.190 182.545 94.445 182.875 ;
        RECT 94.670 182.545 94.865 182.875 ;
        RECT 88.715 181.405 90.745 181.575 ;
        RECT 92.005 181.405 92.275 182.310 ;
        RECT 92.460 182.165 93.125 182.335 ;
        RECT 92.955 181.405 93.125 182.165 ;
        RECT 93.850 181.405 94.185 182.375 ;
        RECT 94.695 181.575 94.865 182.545 ;
        RECT 95.035 181.915 95.205 183.045 ;
        RECT 95.375 182.255 95.545 183.055 ;
        RECT 95.750 182.765 96.025 183.615 ;
        RECT 95.745 182.595 96.025 182.765 ;
        RECT 95.750 182.455 96.025 182.595 ;
        RECT 96.195 182.255 96.385 183.615 ;
        RECT 97.295 182.975 97.540 183.580 ;
        RECT 97.990 183.045 98.245 183.615 ;
        RECT 99.170 183.250 99.700 183.615 ;
        RECT 99.890 183.445 100.165 183.615 ;
        RECT 99.885 183.275 100.165 183.445 ;
        RECT 99.170 183.215 99.345 183.250 ;
        RECT 98.415 183.045 99.345 183.215 ;
        RECT 96.585 182.805 97.815 182.975 ;
        RECT 95.375 182.085 96.385 182.255 ;
        RECT 96.555 182.240 97.305 182.430 ;
        RECT 95.035 181.745 96.160 181.915 ;
        RECT 96.555 181.575 96.725 182.240 ;
        RECT 97.475 181.995 97.815 182.805 ;
        RECT 97.300 181.585 97.815 181.995 ;
        RECT 97.990 182.375 98.160 183.045 ;
        RECT 98.415 182.875 98.585 183.045 ;
        RECT 98.330 182.545 98.585 182.875 ;
        RECT 98.810 182.545 99.005 182.875 ;
        RECT 94.695 181.405 96.725 181.575 ;
        RECT 97.990 181.405 98.325 182.375 ;
        RECT 98.835 181.575 99.005 182.545 ;
        RECT 99.175 181.915 99.345 183.045 ;
        RECT 99.515 182.255 99.685 183.055 ;
        RECT 99.890 182.455 100.165 183.275 ;
        RECT 100.335 182.255 100.525 183.615 ;
        RECT 101.435 182.975 101.680 183.580 ;
        RECT 103.095 183.135 103.265 183.615 ;
        RECT 103.935 183.135 104.105 183.615 ;
        RECT 104.775 183.135 104.945 183.615 ;
        RECT 105.535 183.135 105.865 183.615 ;
        RECT 100.725 182.805 101.955 182.975 ;
        RECT 99.515 182.085 100.525 182.255 ;
        RECT 100.695 182.240 101.445 182.430 ;
        RECT 99.175 181.745 100.300 181.915 ;
        RECT 100.695 181.575 100.865 182.240 ;
        RECT 101.615 181.995 101.955 182.805 ;
        RECT 101.440 181.585 101.955 181.995 ;
        RECT 103.095 182.965 104.945 183.135 ;
        RECT 105.115 182.965 105.865 183.135 ;
        RECT 106.730 183.045 106.985 183.615 ;
        RECT 107.910 183.250 108.440 183.615 ;
        RECT 107.910 183.215 108.085 183.250 ;
        RECT 107.155 183.045 108.085 183.215 ;
        RECT 103.095 182.425 104.430 182.965 ;
        RECT 105.115 182.795 105.285 182.965 ;
        RECT 104.815 182.625 105.285 182.795 ;
        RECT 103.095 182.255 104.945 182.425 ;
        RECT 98.835 181.405 100.865 181.575 ;
        RECT 103.095 181.405 103.265 182.255 ;
        RECT 103.935 181.405 104.105 182.255 ;
        RECT 104.775 181.405 104.945 182.255 ;
        RECT 105.115 182.385 105.285 182.625 ;
        RECT 105.455 182.555 106.360 182.795 ;
        RECT 105.115 182.215 105.865 182.385 ;
        RECT 105.535 181.405 105.865 182.215 ;
        RECT 106.730 182.375 106.900 183.045 ;
        RECT 107.155 182.875 107.325 183.045 ;
        RECT 107.070 182.545 107.325 182.875 ;
        RECT 107.550 182.545 107.745 182.875 ;
        RECT 106.730 181.405 107.065 182.375 ;
        RECT 107.575 181.575 107.745 182.545 ;
        RECT 107.915 181.915 108.085 183.045 ;
        RECT 108.255 182.255 108.425 183.055 ;
        RECT 108.630 182.765 108.905 183.615 ;
        RECT 108.625 182.595 108.905 182.765 ;
        RECT 108.630 182.455 108.905 182.595 ;
        RECT 109.075 182.255 109.265 183.615 ;
        RECT 110.175 182.975 110.420 183.580 ;
        RECT 110.955 183.135 111.125 183.615 ;
        RECT 109.465 182.805 110.695 182.975 ;
        RECT 110.955 182.965 111.590 183.135 ;
        RECT 108.255 182.085 109.265 182.255 ;
        RECT 109.435 182.240 110.185 182.430 ;
        RECT 107.915 181.745 109.040 181.915 ;
        RECT 109.435 181.575 109.605 182.240 ;
        RECT 110.355 181.995 110.695 182.805 ;
        RECT 111.420 182.795 111.590 182.965 ;
        RECT 110.870 182.555 111.250 182.795 ;
        RECT 111.420 182.625 111.920 182.795 ;
        RECT 111.420 182.385 111.590 182.625 ;
        RECT 110.180 181.585 110.695 181.995 ;
        RECT 110.875 182.215 111.590 182.385 ;
        RECT 107.575 181.405 109.605 181.575 ;
        RECT 110.875 181.405 111.205 182.215 ;
        RECT 49.685 179.910 50.025 180.895 ;
        RECT 51.850 180.465 52.175 180.895 ;
        RECT 50.195 180.295 52.175 180.465 ;
        RECT 49.685 179.255 49.940 179.910 ;
        RECT 50.195 179.755 50.460 180.295 ;
        RECT 50.675 179.955 51.300 180.125 ;
        RECT 50.110 179.425 50.460 179.755 ;
        RECT 50.630 179.425 50.960 179.755 ;
        RECT 51.130 179.255 51.300 179.955 ;
        RECT 49.685 178.880 50.045 179.255 ;
        RECT 50.760 179.085 51.300 179.255 ;
        RECT 51.470 179.885 52.175 180.295 ;
        RECT 53.805 179.915 54.135 180.895 ;
        RECT 63.030 179.925 63.365 180.895 ;
        RECT 63.875 180.725 65.905 180.895 ;
        RECT 50.760 178.880 50.930 179.085 ;
        RECT 49.745 178.855 49.915 178.880 ;
        RECT 51.470 178.685 51.640 179.885 ;
        RECT 51.810 179.505 52.380 179.715 ;
        RECT 52.550 179.505 53.195 179.715 ;
        RECT 51.870 179.165 53.040 179.335 ;
        RECT 51.870 178.685 52.200 179.165 ;
        RECT 52.710 178.700 53.040 179.165 ;
        RECT 53.805 179.315 54.055 179.915 ;
        RECT 54.225 179.505 54.555 179.755 ;
        RECT 53.805 178.685 54.135 179.315 ;
        RECT 63.030 179.255 63.200 179.925 ;
        RECT 63.875 179.755 64.045 180.725 ;
        RECT 63.370 179.425 63.625 179.755 ;
        RECT 63.850 179.425 64.045 179.755 ;
        RECT 64.215 180.385 65.340 180.555 ;
        RECT 63.455 179.255 63.625 179.425 ;
        RECT 64.215 179.255 64.385 180.385 ;
        RECT 63.030 178.685 63.285 179.255 ;
        RECT 63.455 179.085 64.385 179.255 ;
        RECT 64.555 180.045 65.565 180.215 ;
        RECT 64.555 179.245 64.725 180.045 ;
        RECT 64.930 179.705 65.205 179.845 ;
        RECT 64.925 179.535 65.205 179.705 ;
        RECT 64.210 179.050 64.385 179.085 ;
        RECT 64.210 178.685 64.740 179.050 ;
        RECT 64.930 178.685 65.205 179.535 ;
        RECT 65.375 178.685 65.565 180.045 ;
        RECT 65.735 180.060 65.905 180.725 ;
        RECT 66.480 180.305 66.995 180.715 ;
        RECT 65.735 179.870 66.485 180.060 ;
        RECT 66.655 179.495 66.995 180.305 ;
        RECT 65.765 179.325 66.995 179.495 ;
        RECT 68.085 179.990 68.355 180.895 ;
        RECT 69.035 180.135 69.215 180.895 ;
        RECT 75.495 180.460 75.680 180.865 ;
        RECT 66.475 178.720 66.720 179.325 ;
        RECT 68.085 179.190 68.265 179.990 ;
        RECT 68.540 179.965 69.215 180.135 ;
        RECT 75.015 180.285 75.680 180.460 ;
        RECT 68.540 179.820 68.710 179.965 ;
        RECT 68.435 179.490 68.710 179.820 ;
        RECT 68.540 179.235 68.710 179.490 ;
        RECT 68.935 179.415 69.275 179.785 ;
        RECT 71.325 179.505 72.955 179.755 ;
        RECT 75.015 179.255 75.355 180.285 ;
        RECT 76.385 180.095 76.655 180.865 ;
        RECT 89.875 180.725 91.905 180.895 ;
        RECT 75.525 179.925 76.655 180.095 ;
        RECT 75.525 179.425 75.775 179.925 ;
        RECT 68.085 178.685 68.345 179.190 ;
        RECT 68.540 179.065 69.205 179.235 ;
        RECT 75.015 179.085 75.700 179.255 ;
        RECT 75.955 179.175 76.315 179.755 ;
        RECT 69.035 178.685 69.205 179.065 ;
        RECT 75.495 178.685 75.700 179.085 ;
        RECT 76.485 179.015 76.655 179.925 ;
        RECT 88.785 180.305 89.300 180.715 ;
        RECT 88.785 179.495 89.125 180.305 ;
        RECT 89.875 180.060 90.045 180.725 ;
        RECT 90.440 180.385 91.565 180.555 ;
        RECT 89.295 179.870 90.045 180.060 ;
        RECT 90.215 180.045 91.225 180.215 ;
        RECT 88.785 179.325 90.015 179.495 ;
        RECT 76.395 178.685 76.655 179.015 ;
        RECT 89.060 178.720 89.305 179.325 ;
        RECT 90.215 178.685 90.405 180.045 ;
        RECT 90.575 179.025 90.850 179.845 ;
        RECT 91.055 179.245 91.225 180.045 ;
        RECT 91.395 179.255 91.565 180.385 ;
        RECT 91.735 179.755 91.905 180.725 ;
        RECT 92.415 179.925 92.750 180.895 ;
        RECT 93.005 180.135 93.185 180.895 ;
        RECT 93.005 179.965 93.680 180.135 ;
        RECT 93.865 179.990 94.135 180.895 ;
        RECT 91.735 179.425 91.930 179.755 ;
        RECT 92.155 179.425 92.410 179.755 ;
        RECT 92.155 179.255 92.325 179.425 ;
        RECT 92.580 179.255 92.750 179.925 ;
        RECT 93.510 179.820 93.680 179.965 ;
        RECT 92.945 179.415 93.285 179.785 ;
        RECT 93.510 179.490 93.785 179.820 ;
        RECT 91.395 179.085 92.325 179.255 ;
        RECT 91.395 179.050 91.570 179.085 ;
        RECT 90.575 178.855 90.855 179.025 ;
        RECT 90.575 178.685 90.850 178.855 ;
        RECT 91.040 178.685 91.570 179.050 ;
        RECT 92.495 178.685 92.750 179.255 ;
        RECT 93.510 179.235 93.680 179.490 ;
        RECT 93.015 179.065 93.680 179.235 ;
        RECT 93.955 179.190 94.135 179.990 ;
        RECT 93.015 178.685 93.185 179.065 ;
        RECT 93.875 178.685 94.135 179.190 ;
        RECT 95.665 179.990 95.920 180.895 ;
        RECT 96.635 180.135 96.805 180.895 ;
        RECT 95.665 179.260 95.835 179.990 ;
        RECT 96.090 179.965 96.805 180.135 ;
        RECT 97.065 179.990 97.335 180.895 ;
        RECT 98.015 180.135 98.185 180.895 ;
        RECT 96.090 179.755 96.260 179.965 ;
        RECT 96.005 179.425 96.260 179.755 ;
        RECT 95.665 178.685 95.920 179.260 ;
        RECT 96.090 179.235 96.260 179.425 ;
        RECT 96.540 179.415 96.895 179.785 ;
        RECT 96.090 179.065 96.805 179.235 ;
        RECT 96.635 178.685 96.805 179.065 ;
        RECT 97.065 179.190 97.235 179.990 ;
        RECT 97.520 179.965 98.185 180.135 ;
        RECT 98.445 179.990 98.715 180.895 ;
        RECT 99.395 180.135 99.565 180.895 ;
        RECT 97.520 179.820 97.690 179.965 ;
        RECT 97.405 179.490 97.690 179.820 ;
        RECT 97.520 179.235 97.690 179.490 ;
        RECT 97.065 178.685 97.325 179.190 ;
        RECT 97.520 179.065 98.185 179.235 ;
        RECT 98.015 178.685 98.185 179.065 ;
        RECT 98.445 179.190 98.615 179.990 ;
        RECT 98.900 179.965 99.565 180.135 ;
        RECT 98.900 179.820 99.070 179.965 ;
        RECT 98.785 179.490 99.070 179.820 ;
        RECT 98.900 179.235 99.070 179.490 ;
        RECT 100.290 179.925 100.625 180.895 ;
        RECT 101.135 180.725 103.165 180.895 ;
        RECT 100.290 179.255 100.460 179.925 ;
        RECT 101.135 179.755 101.305 180.725 ;
        RECT 100.630 179.425 100.885 179.755 ;
        RECT 101.110 179.425 101.305 179.755 ;
        RECT 101.475 180.385 102.600 180.555 ;
        RECT 100.715 179.255 100.885 179.425 ;
        RECT 101.475 179.255 101.645 180.385 ;
        RECT 98.445 178.685 98.705 179.190 ;
        RECT 98.900 179.065 99.565 179.235 ;
        RECT 99.395 178.685 99.565 179.065 ;
        RECT 100.290 178.685 100.545 179.255 ;
        RECT 100.715 179.085 101.645 179.255 ;
        RECT 101.815 180.045 102.825 180.215 ;
        RECT 101.815 179.245 101.985 180.045 ;
        RECT 102.190 179.365 102.465 179.845 ;
        RECT 102.185 179.195 102.465 179.365 ;
        RECT 101.470 179.050 101.645 179.085 ;
        RECT 101.470 178.685 102.000 179.050 ;
        RECT 102.190 178.685 102.465 179.195 ;
        RECT 102.635 178.685 102.825 180.045 ;
        RECT 102.995 180.060 103.165 180.725 ;
        RECT 103.740 180.305 104.255 180.715 ;
        RECT 102.995 179.870 103.745 180.060 ;
        RECT 103.915 179.495 104.255 180.305 ;
        RECT 103.025 179.325 104.255 179.495 ;
        RECT 104.425 179.990 104.695 180.895 ;
        RECT 105.375 180.135 105.555 180.895 ;
        RECT 103.735 178.720 103.980 179.325 ;
        RECT 104.425 179.190 104.605 179.990 ;
        RECT 104.880 179.965 105.555 180.135 ;
        RECT 106.725 180.095 106.995 180.865 ;
        RECT 107.700 180.460 107.885 180.865 ;
        RECT 109.025 180.470 109.460 180.895 ;
        RECT 107.700 180.285 108.365 180.460 ;
        RECT 109.025 180.300 110.015 180.470 ;
        RECT 104.880 179.820 105.050 179.965 ;
        RECT 104.775 179.490 105.050 179.820 ;
        RECT 104.880 179.235 105.050 179.490 ;
        RECT 106.725 179.925 107.855 180.095 ;
        RECT 104.425 178.685 104.685 179.190 ;
        RECT 104.880 179.065 105.545 179.235 ;
        RECT 105.375 178.685 105.545 179.065 ;
        RECT 106.725 179.015 106.895 179.925 ;
        RECT 107.065 179.175 107.425 179.755 ;
        RECT 107.605 179.425 107.855 179.925 ;
        RECT 108.025 179.255 108.365 180.285 ;
        RECT 109.025 179.425 109.510 180.130 ;
        RECT 109.680 179.755 110.015 180.300 ;
        RECT 110.185 180.105 110.610 180.895 ;
        RECT 110.780 180.470 111.055 180.895 ;
        RECT 110.780 180.275 111.610 180.470 ;
        RECT 110.185 179.925 111.090 180.105 ;
        RECT 109.680 179.425 110.090 179.755 ;
        RECT 110.260 179.425 111.090 179.925 ;
        RECT 111.260 179.755 111.610 180.275 ;
        RECT 111.780 180.105 112.025 180.895 ;
        RECT 112.215 180.470 112.470 180.895 ;
        RECT 112.215 180.275 113.025 180.470 ;
        RECT 111.780 179.925 112.505 180.105 ;
        RECT 111.260 179.425 111.685 179.755 ;
        RECT 111.855 179.425 112.505 179.925 ;
        RECT 112.675 179.755 113.025 180.275 ;
        RECT 113.195 179.925 113.455 180.895 ;
        RECT 112.675 179.425 113.100 179.755 ;
        RECT 109.680 179.255 110.015 179.425 ;
        RECT 110.260 179.255 110.610 179.425 ;
        RECT 111.260 179.255 111.610 179.425 ;
        RECT 111.855 179.255 112.025 179.425 ;
        RECT 112.675 179.255 113.025 179.425 ;
        RECT 113.270 179.255 113.455 179.925 ;
        RECT 107.680 179.085 108.365 179.255 ;
        RECT 109.025 179.085 110.015 179.255 ;
        RECT 106.725 178.685 106.985 179.015 ;
        RECT 107.680 178.685 107.885 179.085 ;
        RECT 109.025 178.685 109.460 179.085 ;
        RECT 110.185 178.685 110.610 179.255 ;
        RECT 110.800 179.085 111.610 179.255 ;
        RECT 110.800 178.685 111.055 179.085 ;
        RECT 111.780 178.685 112.025 179.255 ;
        RECT 112.215 179.085 113.025 179.255 ;
        RECT 112.215 178.685 112.470 179.085 ;
        RECT 113.195 178.685 113.455 179.255 ;
        RECT 49.685 177.400 50.025 178.175 ;
        RECT 50.605 177.910 50.965 178.175 ;
        RECT 50.605 177.905 50.960 177.910 ;
        RECT 50.605 177.895 50.955 177.905 ;
        RECT 50.605 177.890 50.950 177.895 ;
        RECT 50.605 177.880 50.945 177.890 ;
        RECT 50.605 177.875 50.940 177.880 ;
        RECT 50.605 177.865 50.930 177.875 ;
        RECT 50.605 177.855 50.920 177.865 ;
        RECT 50.605 177.715 50.905 177.855 ;
        RECT 50.195 177.525 50.905 177.715 ;
        RECT 51.095 177.715 51.425 177.795 ;
        RECT 51.935 177.715 52.275 178.175 ;
        RECT 51.095 177.525 52.275 177.715 ;
        RECT 58.430 177.605 58.685 178.175 ;
        RECT 59.610 177.810 60.140 178.175 ;
        RECT 60.330 178.005 60.605 178.175 ;
        RECT 60.325 177.835 60.605 178.005 ;
        RECT 59.610 177.775 59.785 177.810 ;
        RECT 58.855 177.605 59.785 177.775 ;
        RECT 49.685 175.965 49.965 177.400 ;
        RECT 50.195 176.955 50.480 177.525 ;
        RECT 50.665 177.125 51.135 177.355 ;
        RECT 51.305 177.335 51.635 177.355 ;
        RECT 51.305 177.155 51.755 177.335 ;
        RECT 51.945 177.155 52.275 177.355 ;
        RECT 50.195 176.740 51.345 176.955 ;
        RECT 51.015 175.965 51.345 176.740 ;
        RECT 51.540 176.040 51.755 177.155 ;
        RECT 52.045 176.815 52.275 177.155 ;
        RECT 58.430 176.935 58.600 177.605 ;
        RECT 58.855 177.435 59.025 177.605 ;
        RECT 58.770 177.105 59.025 177.435 ;
        RECT 59.250 177.105 59.445 177.435 ;
        RECT 58.430 175.965 58.765 176.935 ;
        RECT 59.275 176.135 59.445 177.105 ;
        RECT 59.615 176.475 59.785 177.605 ;
        RECT 59.955 176.815 60.125 177.615 ;
        RECT 60.330 177.015 60.605 177.835 ;
        RECT 60.775 176.815 60.965 178.175 ;
        RECT 61.875 177.535 62.120 178.140 ;
        RECT 62.565 177.845 62.865 178.175 ;
        RECT 61.165 177.365 62.395 177.535 ;
        RECT 59.955 176.645 60.965 176.815 ;
        RECT 61.135 176.800 61.885 176.990 ;
        RECT 59.615 176.305 60.740 176.475 ;
        RECT 61.135 176.135 61.305 176.800 ;
        RECT 62.055 176.555 62.395 177.365 ;
        RECT 61.880 176.145 62.395 176.555 ;
        RECT 62.565 176.935 62.735 177.845 ;
        RECT 63.490 177.695 63.785 178.085 ;
        RECT 64.385 177.695 64.645 178.085 ;
        RECT 68.195 177.965 69.365 178.175 ;
        RECT 68.195 177.945 68.525 177.965 ;
        RECT 62.905 177.105 63.255 177.675 ;
        RECT 63.490 177.525 65.140 177.695 ;
        RECT 63.425 177.185 64.565 177.355 ;
        RECT 63.425 176.935 63.595 177.185 ;
        RECT 64.735 177.015 65.140 177.525 ;
        RECT 62.565 176.765 63.595 176.935 ;
        RECT 64.385 176.845 65.140 177.015 ;
        RECT 68.085 177.525 68.945 177.775 ;
        RECT 69.115 177.715 69.365 177.965 ;
        RECT 69.875 177.715 70.215 178.175 ;
        RECT 69.115 177.545 70.215 177.715 ;
        RECT 75.910 177.605 76.165 178.175 ;
        RECT 77.090 177.810 77.620 178.175 ;
        RECT 77.090 177.775 77.265 177.810 ;
        RECT 76.335 177.605 77.265 177.775 ;
        RECT 68.085 176.935 68.365 177.525 ;
        RECT 68.535 177.105 69.285 177.355 ;
        RECT 75.910 176.935 76.080 177.605 ;
        RECT 76.335 177.435 76.505 177.605 ;
        RECT 76.250 177.105 76.505 177.435 ;
        RECT 76.730 177.105 76.925 177.435 ;
        RECT 59.275 175.965 61.305 176.135 ;
        RECT 62.565 175.965 62.875 176.765 ;
        RECT 64.385 176.595 64.645 176.845 ;
        RECT 68.085 176.765 69.785 176.935 ;
        RECT 63.525 176.425 64.645 176.595 ;
        RECT 63.525 175.965 63.785 176.425 ;
        RECT 64.385 175.965 64.645 176.425 ;
        RECT 68.615 175.965 68.945 176.765 ;
        RECT 69.455 175.965 69.785 176.765 ;
        RECT 75.910 175.965 76.245 176.935 ;
        RECT 76.755 176.135 76.925 177.105 ;
        RECT 77.095 176.475 77.265 177.605 ;
        RECT 77.435 176.815 77.605 177.615 ;
        RECT 77.810 177.325 78.085 178.175 ;
        RECT 77.805 177.155 78.085 177.325 ;
        RECT 77.810 177.015 78.085 177.155 ;
        RECT 78.255 176.815 78.445 178.175 ;
        RECT 79.355 177.535 79.600 178.140 ;
        RECT 78.645 177.365 79.875 177.535 ;
        RECT 77.435 176.645 78.445 176.815 ;
        RECT 78.615 176.800 79.365 176.990 ;
        RECT 77.095 176.305 78.220 176.475 ;
        RECT 78.615 176.135 78.785 176.800 ;
        RECT 79.535 176.555 79.875 177.365 ;
        RECT 79.360 176.145 79.875 176.555 ;
        RECT 76.755 175.965 78.785 176.135 ;
        RECT 80.045 175.965 80.305 178.175 ;
        RECT 80.895 178.005 81.890 178.175 ;
        RECT 82.420 178.015 82.590 178.175 ;
        RECT 80.895 177.715 81.065 178.005 ;
        RECT 81.720 177.845 81.890 178.005 ;
        RECT 82.060 177.845 82.590 178.015 ;
        RECT 80.495 177.545 81.065 177.715 ;
        RECT 81.235 177.665 81.410 177.835 ;
        RECT 80.495 176.765 80.665 177.545 ;
        RECT 81.235 177.505 81.650 177.665 ;
        RECT 81.240 177.495 81.650 177.505 ;
        RECT 80.975 177.155 81.430 177.325 ;
        RECT 80.495 176.595 81.145 176.765 ;
        RECT 82.060 176.675 82.230 177.845 ;
        RECT 82.935 177.775 83.110 178.105 ;
        RECT 82.400 177.495 82.640 177.665 ;
        RECT 80.975 176.135 81.145 176.595 ;
        RECT 81.445 176.445 82.230 176.675 ;
        RECT 81.445 176.305 81.775 176.445 ;
        RECT 82.470 176.295 82.640 177.495 ;
        RECT 82.935 177.325 83.105 177.775 ;
        RECT 83.880 177.715 84.125 178.135 ;
        RECT 84.640 178.005 86.240 178.175 ;
        RECT 84.640 177.965 84.995 178.005 ;
        RECT 85.230 177.715 85.400 177.835 ;
        RECT 83.880 177.545 85.400 177.715 ;
        RECT 85.230 177.505 85.400 177.545 ;
        RECT 85.570 177.585 85.900 177.835 ;
        RECT 86.070 177.635 86.240 178.005 ;
        RECT 87.530 178.005 88.605 178.175 ;
        RECT 85.570 177.510 85.885 177.585 ;
        RECT 82.815 177.155 83.105 177.325 ;
        RECT 81.930 176.135 82.260 176.175 ;
        RECT 80.975 175.965 82.260 176.135 ;
        RECT 82.430 175.965 82.640 176.295 ;
        RECT 82.935 176.295 83.105 177.155 ;
        RECT 83.275 176.755 83.565 177.435 ;
        RECT 84.040 176.755 84.370 177.375 ;
        RECT 84.575 177.325 84.820 177.375 ;
        RECT 85.215 177.325 85.545 177.335 ;
        RECT 84.575 177.155 84.875 177.325 ;
        RECT 85.160 177.165 85.545 177.325 ;
        RECT 85.160 177.155 85.330 177.165 ;
        RECT 84.575 176.755 84.820 177.155 ;
        RECT 85.715 176.985 85.885 177.510 ;
        RECT 85.125 176.815 85.885 176.985 ;
        RECT 83.890 176.345 84.955 176.515 ;
        RECT 82.935 175.965 83.120 176.295 ;
        RECT 83.890 175.965 84.060 176.345 ;
        RECT 84.785 176.135 84.955 176.345 ;
        RECT 85.125 176.305 85.455 176.815 ;
        RECT 85.625 176.135 85.795 176.645 ;
        RECT 86.055 176.435 86.355 177.435 ;
        RECT 87.000 177.325 87.360 178.000 ;
        RECT 87.530 177.670 87.700 178.005 ;
        RECT 87.870 177.665 88.210 177.835 ;
        RECT 87.920 177.495 88.210 177.665 ;
        RECT 88.435 177.795 88.605 178.005 ;
        RECT 89.275 177.795 89.445 178.170 ;
        RECT 88.435 177.625 89.445 177.795 ;
        RECT 89.705 177.885 90.265 178.175 ;
        RECT 87.000 177.145 87.540 177.325 ;
        RECT 87.000 177.035 87.360 177.145 ;
        RECT 86.555 176.805 87.360 177.035 ;
        RECT 88.040 176.975 88.210 177.495 ;
        RECT 87.575 176.805 88.210 176.975 ;
        RECT 88.380 176.815 88.815 177.435 ;
        RECT 89.125 176.985 89.470 177.435 ;
        RECT 89.125 176.815 89.475 176.985 ;
        RECT 84.785 175.965 85.795 176.135 ;
        RECT 86.555 175.965 86.905 176.805 ;
        RECT 87.075 176.135 87.245 176.635 ;
        RECT 87.575 176.475 87.745 176.805 ;
        RECT 87.415 176.305 87.745 176.475 ;
        RECT 87.915 176.465 89.445 176.635 ;
        RECT 87.915 176.305 88.085 176.465 ;
        RECT 88.435 176.135 88.605 176.295 ;
        RECT 87.075 175.965 88.605 176.135 ;
        RECT 89.275 175.965 89.445 176.465 ;
        RECT 89.705 176.515 89.955 177.885 ;
        RECT 91.305 177.715 91.635 178.075 ;
        RECT 90.245 177.525 91.635 177.715 ;
        RECT 93.850 177.605 94.105 178.175 ;
        RECT 95.030 177.810 95.560 178.175 ;
        RECT 95.030 177.775 95.205 177.810 ;
        RECT 94.275 177.605 95.205 177.775 ;
        RECT 90.245 177.435 90.415 177.525 ;
        RECT 90.125 177.105 90.415 177.435 ;
        RECT 90.585 177.105 90.925 177.355 ;
        RECT 90.245 176.855 90.415 177.105 ;
        RECT 93.850 176.935 94.020 177.605 ;
        RECT 94.275 177.435 94.445 177.605 ;
        RECT 94.190 177.105 94.445 177.435 ;
        RECT 94.670 177.105 94.865 177.435 ;
        RECT 90.245 176.685 91.185 176.855 ;
        RECT 89.705 175.965 90.165 176.515 ;
        RECT 90.885 176.135 91.185 176.685 ;
        RECT 93.850 175.965 94.185 176.935 ;
        RECT 94.695 176.135 94.865 177.105 ;
        RECT 95.035 176.475 95.205 177.605 ;
        RECT 95.375 176.815 95.545 177.615 ;
        RECT 95.750 177.325 96.025 178.175 ;
        RECT 95.745 177.155 96.025 177.325 ;
        RECT 95.750 177.015 96.025 177.155 ;
        RECT 96.195 176.815 96.385 178.175 ;
        RECT 97.295 177.535 97.540 178.140 ;
        RECT 98.675 177.695 99.005 178.175 ;
        RECT 99.595 177.695 99.765 178.175 ;
        RECT 100.435 177.695 100.605 178.175 ;
        RECT 101.275 177.695 101.445 178.175 ;
        RECT 96.585 177.365 97.815 177.535 ;
        RECT 98.675 177.525 99.425 177.695 ;
        RECT 99.595 177.525 101.445 177.695 ;
        RECT 95.375 176.645 96.385 176.815 ;
        RECT 96.555 176.800 97.305 176.990 ;
        RECT 95.035 176.305 96.160 176.475 ;
        RECT 96.555 176.135 96.725 176.800 ;
        RECT 97.475 176.555 97.815 177.365 ;
        RECT 99.255 177.355 99.425 177.525 ;
        RECT 98.180 177.115 99.085 177.355 ;
        RECT 99.255 177.185 99.725 177.355 ;
        RECT 99.255 176.945 99.425 177.185 ;
        RECT 100.110 176.985 101.445 177.525 ;
        RECT 97.300 176.145 97.815 176.555 ;
        RECT 98.675 176.775 99.425 176.945 ;
        RECT 99.595 176.815 101.445 176.985 ;
        RECT 94.695 175.965 96.725 176.135 ;
        RECT 98.675 175.965 99.005 176.775 ;
        RECT 99.595 175.965 99.765 176.815 ;
        RECT 100.435 175.965 100.605 176.815 ;
        RECT 101.275 175.965 101.445 176.815 ;
        RECT 103.050 177.605 103.305 178.175 ;
        RECT 104.230 177.810 104.760 178.175 ;
        RECT 104.230 177.775 104.405 177.810 ;
        RECT 103.475 177.605 104.405 177.775 ;
        RECT 103.050 176.935 103.220 177.605 ;
        RECT 103.475 177.435 103.645 177.605 ;
        RECT 103.390 177.105 103.645 177.435 ;
        RECT 103.870 177.105 104.065 177.435 ;
        RECT 103.050 175.965 103.385 176.935 ;
        RECT 103.895 176.135 104.065 177.105 ;
        RECT 104.235 176.475 104.405 177.605 ;
        RECT 104.575 176.815 104.745 177.615 ;
        RECT 104.950 177.325 105.225 178.175 ;
        RECT 104.945 177.155 105.225 177.325 ;
        RECT 104.950 177.015 105.225 177.155 ;
        RECT 105.395 176.815 105.585 178.175 ;
        RECT 106.495 177.535 106.740 178.140 ;
        RECT 108.085 177.600 108.340 178.175 ;
        RECT 109.055 177.795 109.225 178.175 ;
        RECT 108.510 177.625 109.225 177.795 ;
        RECT 110.915 177.695 111.085 178.175 ;
        RECT 111.755 177.695 111.925 178.175 ;
        RECT 112.595 177.695 112.765 178.175 ;
        RECT 113.355 177.695 113.685 178.175 ;
        RECT 105.785 177.365 107.015 177.535 ;
        RECT 104.575 176.645 105.585 176.815 ;
        RECT 105.755 176.800 106.505 176.990 ;
        RECT 104.235 176.305 105.360 176.475 ;
        RECT 105.755 176.135 105.925 176.800 ;
        RECT 106.675 176.555 107.015 177.365 ;
        RECT 106.500 176.145 107.015 176.555 ;
        RECT 108.085 176.870 108.255 177.600 ;
        RECT 108.510 177.435 108.680 177.625 ;
        RECT 108.425 177.105 108.680 177.435 ;
        RECT 108.510 176.895 108.680 177.105 ;
        RECT 110.915 177.525 112.765 177.695 ;
        RECT 112.935 177.525 113.685 177.695 ;
        RECT 110.915 176.985 112.250 177.525 ;
        RECT 112.935 177.355 113.105 177.525 ;
        RECT 112.635 177.185 113.105 177.355 ;
        RECT 103.895 175.965 105.925 176.135 ;
        RECT 108.085 175.965 108.340 176.870 ;
        RECT 108.510 176.725 109.225 176.895 ;
        RECT 109.055 175.965 109.225 176.725 ;
        RECT 110.915 176.815 112.765 176.985 ;
        RECT 110.915 175.965 111.085 176.815 ;
        RECT 111.755 175.965 111.925 176.815 ;
        RECT 112.595 175.965 112.765 176.815 ;
        RECT 112.935 176.945 113.105 177.185 ;
        RECT 113.275 177.115 114.180 177.355 ;
        RECT 112.935 176.775 113.685 176.945 ;
        RECT 113.355 175.965 113.685 176.775 ;
        RECT 49.235 174.945 49.565 175.455 ;
        RECT 50.945 175.115 51.325 175.285 ;
        RECT 51.155 174.945 51.325 175.115 ;
        RECT 55.675 174.945 56.005 175.455 ;
        RECT 57.385 175.115 57.765 175.285 ;
        RECT 57.595 174.945 57.765 175.115 ;
        RECT 48.765 174.775 50.985 174.945 ;
        RECT 48.765 173.815 48.935 174.775 ;
        RECT 49.105 174.435 50.645 174.605 ;
        RECT 49.105 173.985 49.350 174.435 ;
        RECT 49.610 174.065 50.305 174.265 ;
        RECT 50.475 174.235 50.645 174.435 ;
        RECT 50.815 174.575 50.985 174.775 ;
        RECT 51.155 174.745 51.815 174.945 ;
        RECT 50.815 174.405 51.475 174.575 ;
        RECT 50.475 174.065 51.075 174.235 ;
        RECT 51.305 173.985 51.475 174.405 ;
        RECT 50.075 173.815 50.985 173.895 ;
        RECT 51.645 173.815 51.815 174.745 ;
        RECT 48.765 173.270 49.230 173.815 ;
        RECT 50.075 173.725 51.325 173.815 ;
        RECT 50.075 173.245 50.405 173.725 ;
        RECT 50.815 173.645 51.325 173.725 ;
        RECT 51.095 173.245 51.325 173.645 ;
        RECT 51.495 173.335 51.815 173.815 ;
        RECT 55.205 174.775 57.425 174.945 ;
        RECT 55.205 173.815 55.375 174.775 ;
        RECT 55.545 174.435 57.085 174.605 ;
        RECT 55.545 173.985 55.790 174.435 ;
        RECT 56.050 174.065 56.745 174.265 ;
        RECT 56.915 174.235 57.085 174.435 ;
        RECT 57.255 174.575 57.425 174.775 ;
        RECT 57.595 174.745 58.255 174.945 ;
        RECT 57.255 174.405 57.915 174.575 ;
        RECT 56.915 174.065 57.515 174.235 ;
        RECT 57.745 173.985 57.915 174.405 ;
        RECT 56.515 173.815 57.425 173.895 ;
        RECT 58.085 173.815 58.255 174.745 ;
        RECT 55.205 173.270 55.670 173.815 ;
        RECT 56.515 173.725 57.765 173.815 ;
        RECT 56.515 173.245 56.845 173.725 ;
        RECT 57.255 173.645 57.765 173.725 ;
        RECT 57.535 173.245 57.765 173.645 ;
        RECT 57.935 173.335 58.255 173.815 ;
        RECT 58.425 174.905 58.885 175.455 ;
        RECT 63.195 175.285 65.225 175.455 ;
        RECT 58.425 173.535 58.675 174.905 ;
        RECT 59.605 174.735 59.905 175.285 ;
        RECT 58.965 174.565 59.905 174.735 ;
        RECT 62.105 174.865 62.620 175.275 ;
        RECT 58.965 174.315 59.135 174.565 ;
        RECT 58.845 173.985 59.135 174.315 ;
        RECT 59.305 174.065 59.645 174.315 ;
        RECT 58.965 173.895 59.135 173.985 ;
        RECT 62.105 174.055 62.445 174.865 ;
        RECT 63.195 174.620 63.365 175.285 ;
        RECT 63.760 174.945 64.885 175.115 ;
        RECT 62.615 174.430 63.365 174.620 ;
        RECT 63.535 174.605 64.545 174.775 ;
        RECT 58.965 173.705 60.355 173.895 ;
        RECT 62.105 173.885 63.335 174.055 ;
        RECT 58.425 173.245 58.985 173.535 ;
        RECT 60.025 173.345 60.355 173.705 ;
        RECT 62.380 173.280 62.625 173.885 ;
        RECT 63.535 173.245 63.725 174.605 ;
        RECT 63.895 173.925 64.170 174.405 ;
        RECT 63.895 173.755 64.175 173.925 ;
        RECT 64.375 173.805 64.545 174.605 ;
        RECT 64.715 173.815 64.885 174.945 ;
        RECT 65.055 174.315 65.225 175.285 ;
        RECT 65.735 174.485 66.070 175.455 ;
        RECT 65.055 173.985 65.250 174.315 ;
        RECT 65.475 173.985 65.730 174.315 ;
        RECT 65.475 173.815 65.645 173.985 ;
        RECT 65.900 173.815 66.070 174.485 ;
        RECT 63.895 173.245 64.170 173.755 ;
        RECT 64.715 173.645 65.645 173.815 ;
        RECT 64.715 173.610 64.890 173.645 ;
        RECT 64.360 173.245 64.890 173.610 ;
        RECT 65.815 173.245 66.070 173.815 ;
        RECT 66.250 174.485 66.585 175.455 ;
        RECT 67.095 175.285 69.125 175.455 ;
        RECT 66.250 173.815 66.420 174.485 ;
        RECT 67.095 174.315 67.265 175.285 ;
        RECT 66.590 173.985 66.845 174.315 ;
        RECT 67.070 173.985 67.265 174.315 ;
        RECT 67.435 174.945 68.560 175.115 ;
        RECT 66.675 173.815 66.845 173.985 ;
        RECT 67.435 173.815 67.605 174.945 ;
        RECT 66.250 173.245 66.505 173.815 ;
        RECT 66.675 173.645 67.605 173.815 ;
        RECT 67.775 174.605 68.785 174.775 ;
        RECT 67.775 173.805 67.945 174.605 ;
        RECT 67.430 173.610 67.605 173.645 ;
        RECT 67.430 173.245 67.960 173.610 ;
        RECT 68.150 173.585 68.425 174.405 ;
        RECT 68.145 173.415 68.425 173.585 ;
        RECT 68.150 173.245 68.425 173.415 ;
        RECT 68.595 173.245 68.785 174.605 ;
        RECT 68.955 174.620 69.125 175.285 ;
        RECT 69.700 174.865 70.215 175.275 ;
        RECT 68.955 174.430 69.705 174.620 ;
        RECT 69.875 174.055 70.215 174.865 ;
        RECT 70.475 174.955 70.645 175.455 ;
        RECT 71.315 175.285 72.845 175.455 ;
        RECT 71.315 175.125 71.485 175.285 ;
        RECT 71.835 174.955 72.005 175.115 ;
        RECT 70.475 174.785 72.005 174.955 ;
        RECT 72.175 174.945 72.505 175.115 ;
        RECT 72.175 174.615 72.345 174.945 ;
        RECT 72.675 174.785 72.845 175.285 ;
        RECT 73.015 174.615 73.365 175.455 ;
        RECT 74.125 175.285 75.135 175.455 ;
        RECT 70.450 174.265 70.795 174.605 ;
        RECT 70.445 174.095 70.795 174.265 ;
        RECT 68.985 173.885 70.215 174.055 ;
        RECT 70.450 173.985 70.795 174.095 ;
        RECT 71.105 173.985 71.540 174.605 ;
        RECT 71.710 174.445 72.345 174.615 ;
        RECT 71.710 173.925 71.880 174.445 ;
        RECT 72.560 174.385 73.365 174.615 ;
        RECT 72.560 174.275 72.920 174.385 ;
        RECT 72.380 174.095 72.920 174.275 ;
        RECT 69.695 173.280 69.940 173.885 ;
        RECT 70.475 173.625 71.485 173.795 ;
        RECT 70.475 173.250 70.645 173.625 ;
        RECT 71.315 173.415 71.485 173.625 ;
        RECT 71.710 173.755 72.000 173.925 ;
        RECT 71.710 173.585 72.050 173.755 ;
        RECT 72.220 173.415 72.390 173.750 ;
        RECT 72.560 173.420 72.920 174.095 ;
        RECT 73.565 173.985 73.865 174.985 ;
        RECT 74.125 174.775 74.295 175.285 ;
        RECT 74.465 174.605 74.795 175.115 ;
        RECT 74.965 175.075 75.135 175.285 ;
        RECT 75.860 175.075 76.030 175.455 ;
        RECT 76.800 175.125 76.985 175.455 ;
        RECT 74.965 174.905 76.030 175.075 ;
        RECT 74.035 174.435 74.795 174.605 ;
        RECT 74.035 173.910 74.205 174.435 ;
        RECT 75.100 174.265 75.345 174.665 ;
        RECT 74.590 174.255 74.760 174.265 ;
        RECT 74.375 174.095 74.760 174.255 ;
        RECT 75.045 174.095 75.345 174.265 ;
        RECT 74.375 174.085 74.705 174.095 ;
        RECT 75.100 174.045 75.345 174.095 ;
        RECT 75.550 174.045 75.880 174.665 ;
        RECT 76.355 173.985 76.645 174.665 ;
        RECT 76.815 174.265 76.985 175.125 ;
        RECT 77.280 175.125 77.490 175.455 ;
        RECT 77.660 175.285 78.945 175.455 ;
        RECT 77.660 175.245 77.990 175.285 ;
        RECT 76.815 174.095 77.105 174.265 ;
        RECT 74.035 173.835 74.350 173.910 ;
        RECT 71.315 173.245 72.390 173.415 ;
        RECT 73.680 173.415 73.850 173.785 ;
        RECT 74.020 173.585 74.350 173.835 ;
        RECT 74.520 173.875 74.690 173.915 ;
        RECT 74.520 173.705 76.040 173.875 ;
        RECT 74.520 173.585 74.690 173.705 ;
        RECT 74.925 173.415 75.280 173.455 ;
        RECT 73.680 173.245 75.280 173.415 ;
        RECT 75.795 173.285 76.040 173.705 ;
        RECT 76.815 173.645 76.985 174.095 ;
        RECT 77.280 173.925 77.450 175.125 ;
        RECT 78.145 174.975 78.475 175.115 ;
        RECT 77.690 174.745 78.475 174.975 ;
        RECT 78.775 174.825 78.945 175.285 ;
        RECT 77.280 173.755 77.520 173.925 ;
        RECT 76.810 173.315 76.985 173.645 ;
        RECT 77.690 173.575 77.860 174.745 ;
        RECT 78.775 174.655 79.425 174.825 ;
        RECT 78.490 174.095 78.945 174.265 ;
        RECT 78.270 173.915 78.680 173.925 ;
        RECT 78.270 173.755 78.685 173.915 ;
        RECT 79.255 173.875 79.425 174.655 ;
        RECT 78.510 173.585 78.685 173.755 ;
        RECT 78.855 173.705 79.425 173.875 ;
        RECT 77.330 173.405 77.860 173.575 ;
        RECT 78.030 173.415 78.200 173.575 ;
        RECT 78.855 173.415 79.025 173.705 ;
        RECT 77.330 173.245 77.500 173.405 ;
        RECT 78.030 173.245 79.025 173.415 ;
        RECT 79.615 173.245 79.875 175.455 ;
        RECT 82.055 175.285 84.085 175.455 ;
        RECT 80.965 174.865 81.480 175.275 ;
        RECT 80.965 174.055 81.305 174.865 ;
        RECT 82.055 174.620 82.225 175.285 ;
        RECT 82.620 174.945 83.745 175.115 ;
        RECT 81.475 174.430 82.225 174.620 ;
        RECT 82.395 174.605 83.405 174.775 ;
        RECT 80.965 173.885 82.195 174.055 ;
        RECT 81.240 173.280 81.485 173.885 ;
        RECT 82.395 173.245 82.585 174.605 ;
        RECT 82.755 173.925 83.030 174.405 ;
        RECT 82.755 173.755 83.035 173.925 ;
        RECT 83.235 173.805 83.405 174.605 ;
        RECT 83.575 173.815 83.745 174.945 ;
        RECT 83.915 174.315 84.085 175.285 ;
        RECT 84.595 174.485 84.930 175.455 ;
        RECT 83.915 173.985 84.110 174.315 ;
        RECT 84.335 173.985 84.590 174.315 ;
        RECT 84.335 173.815 84.505 173.985 ;
        RECT 84.760 173.815 84.930 174.485 ;
        RECT 82.755 173.245 83.030 173.755 ;
        RECT 83.575 173.645 84.505 173.815 ;
        RECT 83.575 173.610 83.750 173.645 ;
        RECT 83.220 173.245 83.750 173.610 ;
        RECT 84.675 173.245 84.930 173.815 ;
        RECT 85.105 174.550 85.375 175.455 ;
        RECT 86.055 174.695 86.235 175.455 ;
        RECT 89.415 175.285 91.445 175.455 ;
        RECT 85.105 173.750 85.285 174.550 ;
        RECT 85.560 174.525 86.235 174.695 ;
        RECT 88.325 174.865 88.840 175.275 ;
        RECT 85.560 174.380 85.730 174.525 ;
        RECT 85.455 174.050 85.730 174.380 ;
        RECT 85.560 173.795 85.730 174.050 ;
        RECT 85.955 173.975 86.295 174.345 ;
        RECT 88.325 174.055 88.665 174.865 ;
        RECT 89.415 174.620 89.585 175.285 ;
        RECT 89.980 174.945 91.105 175.115 ;
        RECT 88.835 174.430 89.585 174.620 ;
        RECT 89.755 174.605 90.765 174.775 ;
        RECT 88.325 173.885 89.555 174.055 ;
        RECT 85.105 173.245 85.365 173.750 ;
        RECT 85.560 173.625 86.225 173.795 ;
        RECT 86.055 173.245 86.225 173.625 ;
        RECT 88.600 173.280 88.845 173.885 ;
        RECT 89.755 173.245 89.945 174.605 ;
        RECT 90.115 174.265 90.390 174.405 ;
        RECT 90.115 174.095 90.395 174.265 ;
        RECT 90.115 173.245 90.390 174.095 ;
        RECT 90.595 173.805 90.765 174.605 ;
        RECT 90.935 173.815 91.105 174.945 ;
        RECT 91.275 174.315 91.445 175.285 ;
        RECT 91.955 174.485 92.290 175.455 ;
        RECT 93.555 175.285 95.585 175.455 ;
        RECT 91.275 173.985 91.470 174.315 ;
        RECT 91.695 173.985 91.950 174.315 ;
        RECT 91.695 173.815 91.865 173.985 ;
        RECT 92.120 173.815 92.290 174.485 ;
        RECT 92.465 174.865 92.980 175.275 ;
        RECT 92.465 174.055 92.805 174.865 ;
        RECT 93.555 174.620 93.725 175.285 ;
        RECT 94.120 174.945 95.245 175.115 ;
        RECT 92.975 174.430 93.725 174.620 ;
        RECT 93.895 174.605 94.905 174.775 ;
        RECT 92.465 173.885 93.695 174.055 ;
        RECT 90.935 173.645 91.865 173.815 ;
        RECT 90.935 173.610 91.110 173.645 ;
        RECT 90.580 173.245 91.110 173.610 ;
        RECT 92.035 173.245 92.290 173.815 ;
        RECT 92.740 173.280 92.985 173.885 ;
        RECT 93.895 173.245 94.085 174.605 ;
        RECT 94.255 173.585 94.530 174.405 ;
        RECT 94.735 173.805 94.905 174.605 ;
        RECT 95.075 173.815 95.245 174.945 ;
        RECT 95.415 174.315 95.585 175.285 ;
        RECT 96.095 174.485 96.430 175.455 ;
        RECT 95.415 173.985 95.610 174.315 ;
        RECT 95.835 173.985 96.090 174.315 ;
        RECT 95.835 173.815 96.005 173.985 ;
        RECT 96.260 173.815 96.430 174.485 ;
        RECT 95.075 173.645 96.005 173.815 ;
        RECT 95.075 173.610 95.250 173.645 ;
        RECT 94.255 173.415 94.535 173.585 ;
        RECT 94.255 173.245 94.530 173.415 ;
        RECT 94.720 173.245 95.250 173.610 ;
        RECT 96.175 173.245 96.430 173.815 ;
        RECT 97.530 174.485 97.865 175.455 ;
        RECT 98.375 175.285 100.405 175.455 ;
        RECT 97.530 173.815 97.700 174.485 ;
        RECT 98.375 174.315 98.545 175.285 ;
        RECT 97.870 173.985 98.125 174.315 ;
        RECT 98.350 173.985 98.545 174.315 ;
        RECT 98.715 174.945 99.840 175.115 ;
        RECT 97.955 173.815 98.125 173.985 ;
        RECT 98.715 173.815 98.885 174.945 ;
        RECT 97.530 173.245 97.785 173.815 ;
        RECT 97.955 173.645 98.885 173.815 ;
        RECT 99.055 174.605 100.065 174.775 ;
        RECT 99.055 173.805 99.225 174.605 ;
        RECT 99.430 173.925 99.705 174.405 ;
        RECT 99.425 173.755 99.705 173.925 ;
        RECT 98.710 173.610 98.885 173.645 ;
        RECT 98.710 173.245 99.240 173.610 ;
        RECT 99.430 173.245 99.705 173.755 ;
        RECT 99.875 173.245 100.065 174.605 ;
        RECT 100.235 174.620 100.405 175.285 ;
        RECT 100.980 174.865 101.495 175.275 ;
        RECT 100.235 174.430 100.985 174.620 ;
        RECT 101.155 174.055 101.495 174.865 ;
        RECT 100.265 173.885 101.495 174.055 ;
        RECT 101.670 174.485 102.005 175.455 ;
        RECT 102.515 175.285 104.545 175.455 ;
        RECT 100.975 173.280 101.220 173.885 ;
        RECT 101.670 173.815 101.840 174.485 ;
        RECT 102.515 174.315 102.685 175.285 ;
        RECT 102.010 173.985 102.265 174.315 ;
        RECT 102.490 173.985 102.685 174.315 ;
        RECT 102.855 174.945 103.980 175.115 ;
        RECT 102.095 173.815 102.265 173.985 ;
        RECT 102.855 173.815 103.025 174.945 ;
        RECT 101.670 173.245 101.925 173.815 ;
        RECT 102.095 173.645 103.025 173.815 ;
        RECT 103.195 174.605 104.205 174.775 ;
        RECT 103.195 173.805 103.365 174.605 ;
        RECT 103.570 174.265 103.845 174.405 ;
        RECT 103.565 174.095 103.845 174.265 ;
        RECT 102.850 173.610 103.025 173.645 ;
        RECT 102.850 173.245 103.380 173.610 ;
        RECT 103.570 173.245 103.845 174.095 ;
        RECT 104.015 173.245 104.205 174.605 ;
        RECT 104.375 174.620 104.545 175.285 ;
        RECT 105.120 174.865 105.635 175.275 ;
        RECT 104.375 174.430 105.125 174.620 ;
        RECT 105.295 174.055 105.635 174.865 ;
        RECT 104.405 173.885 105.635 174.055 ;
        RECT 106.730 174.485 107.065 175.455 ;
        RECT 107.575 175.285 109.605 175.455 ;
        RECT 105.115 173.280 105.360 173.885 ;
        RECT 106.730 173.815 106.900 174.485 ;
        RECT 107.575 174.315 107.745 175.285 ;
        RECT 107.070 173.985 107.325 174.315 ;
        RECT 107.550 173.985 107.745 174.315 ;
        RECT 107.915 174.945 109.040 175.115 ;
        RECT 107.155 173.815 107.325 173.985 ;
        RECT 107.915 173.815 108.085 174.945 ;
        RECT 106.730 173.245 106.985 173.815 ;
        RECT 107.155 173.645 108.085 173.815 ;
        RECT 108.255 174.605 109.265 174.775 ;
        RECT 108.255 173.805 108.425 174.605 ;
        RECT 108.630 174.265 108.905 174.405 ;
        RECT 108.625 174.095 108.905 174.265 ;
        RECT 107.910 173.610 108.085 173.645 ;
        RECT 107.910 173.245 108.440 173.610 ;
        RECT 108.630 173.245 108.905 174.095 ;
        RECT 109.075 173.245 109.265 174.605 ;
        RECT 109.435 174.620 109.605 175.285 ;
        RECT 110.180 174.865 110.695 175.275 ;
        RECT 109.435 174.430 110.185 174.620 ;
        RECT 110.355 174.055 110.695 174.865 ;
        RECT 109.465 173.885 110.695 174.055 ;
        RECT 112.435 174.605 112.605 175.455 ;
        RECT 113.275 174.605 113.445 175.455 ;
        RECT 114.035 174.645 114.365 175.455 ;
        RECT 112.435 174.435 113.445 174.605 ;
        RECT 113.650 174.475 114.365 174.645 ;
        RECT 112.435 173.895 112.930 174.435 ;
        RECT 113.650 174.235 113.820 174.475 ;
        RECT 113.320 174.065 113.820 174.235 ;
        RECT 113.650 173.895 113.820 174.065 ;
        RECT 110.175 173.280 110.420 173.885 ;
        RECT 112.435 173.725 113.445 173.895 ;
        RECT 113.650 173.725 114.285 173.895 ;
        RECT 112.435 173.245 112.605 173.725 ;
        RECT 113.275 173.245 113.445 173.725 ;
        RECT 114.115 173.245 114.285 173.725 ;
        RECT 56.130 172.165 56.385 172.735 ;
        RECT 57.310 172.370 57.840 172.735 ;
        RECT 57.310 172.335 57.485 172.370 ;
        RECT 56.555 172.165 57.485 172.335 ;
        RECT 56.130 171.495 56.300 172.165 ;
        RECT 56.555 171.995 56.725 172.165 ;
        RECT 56.470 171.665 56.725 171.995 ;
        RECT 56.950 171.665 57.145 171.995 ;
        RECT 56.130 170.525 56.465 171.495 ;
        RECT 56.975 170.695 57.145 171.665 ;
        RECT 57.315 171.035 57.485 172.165 ;
        RECT 57.655 171.375 57.825 172.175 ;
        RECT 58.030 171.885 58.305 172.735 ;
        RECT 58.025 171.715 58.305 171.885 ;
        RECT 58.030 171.575 58.305 171.715 ;
        RECT 58.475 171.375 58.665 172.735 ;
        RECT 59.575 172.095 59.820 172.700 ;
        RECT 62.615 172.335 62.875 172.735 ;
        RECT 64.135 172.350 64.465 172.735 ;
        RECT 64.135 172.335 64.725 172.350 ;
        RECT 62.615 172.165 64.725 172.335 ;
        RECT 58.865 171.925 60.095 172.095 ;
        RECT 57.655 171.205 58.665 171.375 ;
        RECT 58.835 171.360 59.585 171.550 ;
        RECT 57.315 170.865 58.440 171.035 ;
        RECT 58.835 170.695 59.005 171.360 ;
        RECT 59.755 171.115 60.095 171.925 ;
        RECT 59.580 170.705 60.095 171.115 ;
        RECT 62.615 170.865 62.875 172.165 ;
        RECT 63.090 171.665 63.605 171.995 ;
        RECT 63.090 170.865 63.260 171.665 ;
        RECT 63.980 171.375 64.385 171.995 ;
        RECT 64.555 171.495 64.725 172.165 ;
        RECT 64.895 171.665 65.235 172.225 ;
        RECT 65.735 172.165 66.075 172.735 ;
        RECT 68.175 172.355 68.345 172.735 ;
        RECT 68.175 172.185 68.840 172.355 ;
        RECT 69.035 172.230 69.295 172.735 ;
        RECT 65.405 171.665 65.680 171.995 ;
        RECT 65.405 171.495 65.575 171.665 ;
        RECT 65.850 171.495 66.075 172.165 ;
        RECT 68.105 171.635 68.445 172.005 ;
        RECT 68.670 171.930 68.840 172.185 ;
        RECT 64.555 171.325 65.575 171.495 ;
        RECT 64.555 171.175 64.725 171.325 ;
        RECT 64.135 170.910 64.725 171.175 ;
        RECT 63.085 170.695 63.260 170.865 ;
        RECT 65.745 170.830 66.075 171.495 ;
        RECT 68.670 171.600 68.945 171.930 ;
        RECT 68.670 171.455 68.840 171.600 ;
        RECT 56.975 170.525 59.005 170.695 ;
        RECT 63.090 170.530 63.260 170.695 ;
        RECT 65.735 170.525 66.075 170.830 ;
        RECT 68.165 171.285 68.840 171.455 ;
        RECT 69.115 171.430 69.295 172.230 ;
        RECT 68.165 170.525 68.345 171.285 ;
        RECT 69.025 170.525 69.295 171.430 ;
        RECT 80.970 172.165 81.225 172.735 ;
        RECT 82.150 172.370 82.680 172.735 ;
        RECT 82.150 172.335 82.325 172.370 ;
        RECT 81.395 172.165 82.325 172.335 ;
        RECT 80.970 171.495 81.140 172.165 ;
        RECT 81.395 171.995 81.565 172.165 ;
        RECT 81.310 171.665 81.565 171.995 ;
        RECT 81.790 171.665 81.985 171.995 ;
        RECT 80.970 170.525 81.305 171.495 ;
        RECT 81.815 170.695 81.985 171.665 ;
        RECT 82.155 171.035 82.325 172.165 ;
        RECT 82.495 171.375 82.665 172.175 ;
        RECT 82.870 171.885 83.145 172.735 ;
        RECT 82.865 171.715 83.145 171.885 ;
        RECT 82.870 171.575 83.145 171.715 ;
        RECT 83.315 171.375 83.505 172.735 ;
        RECT 84.415 172.095 84.660 172.700 ;
        RECT 86.025 172.330 86.575 172.735 ;
        RECT 87.900 172.330 88.230 172.735 ;
        RECT 89.315 172.500 89.645 172.735 ;
        RECT 86.025 172.275 88.230 172.330 ;
        RECT 89.395 172.275 89.645 172.500 ;
        RECT 90.155 172.275 90.485 172.735 ;
        RECT 97.065 172.330 97.615 172.735 ;
        RECT 98.940 172.330 99.270 172.735 ;
        RECT 100.355 172.500 100.685 172.735 ;
        RECT 97.065 172.275 99.270 172.330 ;
        RECT 100.435 172.275 100.685 172.500 ;
        RECT 101.195 172.275 101.525 172.735 ;
        RECT 104.975 172.355 105.145 172.730 ;
        RECT 105.815 172.565 106.890 172.735 ;
        RECT 105.815 172.355 105.985 172.565 ;
        RECT 86.025 172.105 89.225 172.275 ;
        RECT 83.705 171.925 84.935 172.095 ;
        RECT 82.495 171.205 83.505 171.375 ;
        RECT 83.675 171.360 84.425 171.550 ;
        RECT 82.155 170.865 83.280 171.035 ;
        RECT 83.675 170.695 83.845 171.360 ;
        RECT 84.595 171.115 84.935 171.925 ;
        RECT 84.420 170.705 84.935 171.115 ;
        RECT 86.025 171.535 86.195 172.105 ;
        RECT 86.365 171.705 86.830 171.915 ;
        RECT 81.815 170.525 83.845 170.695 ;
        RECT 86.025 170.525 86.405 171.535 ;
        RECT 86.660 171.075 86.830 171.705 ;
        RECT 87.000 171.355 87.390 171.915 ;
        RECT 87.560 171.445 87.730 172.105 ;
        RECT 89.055 171.915 89.225 172.105 ;
        RECT 89.395 172.085 90.915 172.275 ;
        RECT 87.900 171.665 88.230 171.915 ;
        RECT 88.400 171.745 88.885 171.915 ;
        RECT 87.560 171.245 88.230 171.445 ;
        RECT 86.660 170.905 87.730 171.075 ;
        RECT 87.900 170.935 88.230 171.245 ;
        RECT 87.560 170.765 87.730 170.905 ;
        RECT 88.400 170.865 88.570 171.745 ;
        RECT 89.055 171.705 90.485 171.915 ;
        RECT 90.655 171.535 90.915 172.085 ;
        RECT 88.385 170.765 88.570 170.865 ;
        RECT 87.560 170.595 88.570 170.765 ;
        RECT 89.315 171.365 90.915 171.535 ;
        RECT 97.065 172.105 100.265 172.275 ;
        RECT 97.065 171.535 97.235 172.105 ;
        RECT 97.405 171.705 97.870 171.915 ;
        RECT 89.315 170.525 89.645 171.365 ;
        RECT 90.155 170.525 90.485 171.365 ;
        RECT 97.065 170.525 97.445 171.535 ;
        RECT 97.700 171.075 97.870 171.705 ;
        RECT 98.040 171.355 98.430 171.915 ;
        RECT 98.600 171.445 98.770 172.105 ;
        RECT 100.095 171.915 100.265 172.105 ;
        RECT 100.435 172.085 101.955 172.275 ;
        RECT 104.975 172.185 105.985 172.355 ;
        RECT 106.210 172.225 106.550 172.395 ;
        RECT 106.720 172.230 106.890 172.565 ;
        RECT 108.180 172.565 109.780 172.735 ;
        RECT 98.940 171.665 99.270 171.915 ;
        RECT 99.440 171.745 99.925 171.915 ;
        RECT 98.600 171.245 99.270 171.445 ;
        RECT 97.700 170.905 98.770 171.075 ;
        RECT 98.940 170.935 99.270 171.245 ;
        RECT 98.600 170.765 98.770 170.905 ;
        RECT 99.440 170.865 99.610 171.745 ;
        RECT 100.095 171.705 101.525 171.915 ;
        RECT 101.695 171.535 101.955 172.085 ;
        RECT 106.210 172.055 106.500 172.225 ;
        RECT 104.950 171.885 105.295 171.995 ;
        RECT 104.945 171.715 105.295 171.885 ;
        RECT 99.425 170.765 99.610 170.865 ;
        RECT 98.600 170.595 99.610 170.765 ;
        RECT 100.355 171.365 101.955 171.535 ;
        RECT 104.950 171.375 105.295 171.715 ;
        RECT 105.605 171.375 106.040 171.995 ;
        RECT 106.210 171.535 106.380 172.055 ;
        RECT 107.060 171.885 107.420 172.560 ;
        RECT 108.180 172.195 108.350 172.565 ;
        RECT 109.425 172.525 109.780 172.565 ;
        RECT 108.520 172.145 108.850 172.395 ;
        RECT 108.535 172.070 108.850 172.145 ;
        RECT 109.020 172.275 109.190 172.395 ;
        RECT 110.295 172.275 110.540 172.695 ;
        RECT 111.310 172.335 111.485 172.665 ;
        RECT 111.830 172.575 112.000 172.735 ;
        RECT 111.830 172.405 112.360 172.575 ;
        RECT 112.530 172.565 113.525 172.735 ;
        RECT 112.530 172.405 112.700 172.565 ;
        RECT 109.020 172.105 110.540 172.275 ;
        RECT 106.880 171.705 107.420 171.885 ;
        RECT 107.060 171.595 107.420 171.705 ;
        RECT 106.210 171.365 106.845 171.535 ;
        RECT 107.060 171.365 107.865 171.595 ;
        RECT 100.355 170.525 100.685 171.365 ;
        RECT 101.195 170.525 101.525 171.365 ;
        RECT 104.975 171.025 106.505 171.195 ;
        RECT 104.975 170.525 105.145 171.025 ;
        RECT 106.335 170.865 106.505 171.025 ;
        RECT 106.675 171.035 106.845 171.365 ;
        RECT 106.675 170.865 107.005 171.035 ;
        RECT 105.815 170.695 105.985 170.855 ;
        RECT 107.175 170.695 107.345 171.195 ;
        RECT 105.815 170.525 107.345 170.695 ;
        RECT 107.515 170.525 107.865 171.365 ;
        RECT 108.065 170.995 108.365 171.995 ;
        RECT 108.535 171.545 108.705 172.070 ;
        RECT 109.020 172.065 109.190 172.105 ;
        RECT 108.875 171.885 109.205 171.895 ;
        RECT 109.600 171.885 109.845 171.935 ;
        RECT 108.875 171.725 109.260 171.885 ;
        RECT 109.090 171.715 109.260 171.725 ;
        RECT 109.545 171.715 109.845 171.885 ;
        RECT 108.535 171.375 109.295 171.545 ;
        RECT 108.625 170.695 108.795 171.205 ;
        RECT 108.965 170.865 109.295 171.375 ;
        RECT 109.600 171.315 109.845 171.715 ;
        RECT 110.050 171.315 110.380 171.935 ;
        RECT 110.855 171.315 111.145 171.995 ;
        RECT 111.315 171.885 111.485 172.335 ;
        RECT 111.780 172.055 112.020 172.225 ;
        RECT 111.315 171.715 111.605 171.885 ;
        RECT 109.465 170.905 110.530 171.075 ;
        RECT 109.465 170.695 109.635 170.905 ;
        RECT 108.625 170.525 109.635 170.695 ;
        RECT 110.360 170.525 110.530 170.905 ;
        RECT 111.315 170.855 111.485 171.715 ;
        RECT 111.300 170.525 111.485 170.855 ;
        RECT 111.780 170.855 111.950 172.055 ;
        RECT 112.190 171.235 112.360 172.405 ;
        RECT 113.010 172.225 113.185 172.395 ;
        RECT 112.770 172.065 113.185 172.225 ;
        RECT 113.355 172.275 113.525 172.565 ;
        RECT 113.355 172.105 113.925 172.275 ;
        RECT 112.770 172.055 113.180 172.065 ;
        RECT 112.990 171.715 113.445 171.885 ;
        RECT 113.755 171.325 113.925 172.105 ;
        RECT 112.190 171.005 112.975 171.235 ;
        RECT 112.645 170.865 112.975 171.005 ;
        RECT 113.275 171.155 113.925 171.325 ;
        RECT 111.780 170.525 111.990 170.855 ;
        RECT 112.160 170.695 112.490 170.735 ;
        RECT 113.275 170.695 113.445 171.155 ;
        RECT 112.160 170.525 113.445 170.695 ;
        RECT 114.115 170.525 114.375 172.735 ;
        RECT 61.355 169.845 63.385 170.015 ;
        RECT 60.265 169.425 60.780 169.835 ;
        RECT 60.265 168.615 60.605 169.425 ;
        RECT 61.355 169.180 61.525 169.845 ;
        RECT 61.920 169.505 63.045 169.675 ;
        RECT 60.775 168.990 61.525 169.180 ;
        RECT 61.695 169.165 62.705 169.335 ;
        RECT 60.265 168.445 61.495 168.615 ;
        RECT 60.540 167.840 60.785 168.445 ;
        RECT 61.695 167.805 61.885 169.165 ;
        RECT 62.055 168.145 62.330 168.965 ;
        RECT 62.535 168.365 62.705 169.165 ;
        RECT 62.875 168.375 63.045 169.505 ;
        RECT 63.215 168.875 63.385 169.845 ;
        RECT 63.895 169.045 64.230 170.015 ;
        RECT 63.215 168.545 63.410 168.875 ;
        RECT 63.635 168.545 63.890 168.875 ;
        RECT 63.635 168.375 63.805 168.545 ;
        RECT 64.060 168.375 64.230 169.045 ;
        RECT 62.875 168.205 63.805 168.375 ;
        RECT 62.875 168.170 63.050 168.205 ;
        RECT 62.055 167.975 62.335 168.145 ;
        RECT 62.055 167.805 62.330 167.975 ;
        RECT 62.520 167.805 63.050 168.170 ;
        RECT 63.975 167.805 64.230 168.375 ;
        RECT 67.625 169.555 68.155 170.015 ;
        RECT 69.295 169.555 69.625 170.015 ;
        RECT 67.625 169.385 69.625 169.555 ;
        RECT 67.625 168.375 67.795 169.385 ;
        RECT 67.965 169.045 70.610 169.215 ;
        RECT 70.825 169.045 71.155 170.015 ;
        RECT 67.965 168.545 68.315 169.045 ;
        RECT 69.955 168.965 70.610 169.045 ;
        RECT 68.545 168.545 69.235 168.875 ;
        RECT 69.405 168.545 69.695 168.875 ;
        RECT 70.465 168.625 70.815 168.795 ;
        RECT 70.465 168.375 70.645 168.625 ;
        RECT 70.985 168.455 71.155 169.045 ;
        RECT 67.625 168.205 70.645 168.375 ;
        RECT 67.625 167.830 68.065 168.205 ;
        RECT 69.295 167.805 69.625 168.205 ;
        RECT 70.825 167.805 71.155 168.455 ;
        RECT 71.770 169.045 72.105 170.015 ;
        RECT 72.615 169.845 74.645 170.015 ;
        RECT 71.770 168.375 71.940 169.045 ;
        RECT 72.615 168.875 72.785 169.845 ;
        RECT 72.110 168.545 72.365 168.875 ;
        RECT 72.590 168.545 72.785 168.875 ;
        RECT 72.955 169.505 74.080 169.675 ;
        RECT 72.195 168.375 72.365 168.545 ;
        RECT 72.955 168.375 73.125 169.505 ;
        RECT 71.770 167.805 72.025 168.375 ;
        RECT 72.195 168.205 73.125 168.375 ;
        RECT 73.295 169.165 74.305 169.335 ;
        RECT 73.295 168.365 73.465 169.165 ;
        RECT 73.670 168.825 73.945 168.965 ;
        RECT 73.665 168.655 73.945 168.825 ;
        RECT 72.950 168.170 73.125 168.205 ;
        RECT 72.950 167.805 73.480 168.170 ;
        RECT 73.670 167.805 73.945 168.655 ;
        RECT 74.115 167.805 74.305 169.165 ;
        RECT 74.475 169.180 74.645 169.845 ;
        RECT 75.220 169.425 75.735 169.835 ;
        RECT 74.475 168.990 75.225 169.180 ;
        RECT 75.395 168.615 75.735 169.425 ;
        RECT 81.975 169.515 82.145 170.015 ;
        RECT 82.815 169.845 84.345 170.015 ;
        RECT 82.815 169.685 82.985 169.845 ;
        RECT 83.335 169.515 83.505 169.675 ;
        RECT 81.975 169.345 83.505 169.515 ;
        RECT 83.675 169.505 84.005 169.675 ;
        RECT 83.675 169.175 83.845 169.505 ;
        RECT 84.175 169.345 84.345 169.845 ;
        RECT 84.515 169.175 84.865 170.015 ;
        RECT 85.625 169.845 86.635 170.015 ;
        RECT 81.950 168.825 82.295 169.165 ;
        RECT 81.945 168.655 82.295 168.825 ;
        RECT 74.505 168.445 75.735 168.615 ;
        RECT 81.950 168.545 82.295 168.655 ;
        RECT 82.605 168.545 83.040 169.165 ;
        RECT 83.210 169.005 83.845 169.175 ;
        RECT 83.210 168.485 83.380 169.005 ;
        RECT 84.060 168.945 84.865 169.175 ;
        RECT 84.060 168.835 84.420 168.945 ;
        RECT 83.880 168.655 84.420 168.835 ;
        RECT 75.215 167.840 75.460 168.445 ;
        RECT 81.975 168.185 82.985 168.355 ;
        RECT 81.975 167.810 82.145 168.185 ;
        RECT 82.815 167.975 82.985 168.185 ;
        RECT 83.210 168.315 83.500 168.485 ;
        RECT 83.210 168.145 83.550 168.315 ;
        RECT 83.720 167.975 83.890 168.310 ;
        RECT 84.060 167.980 84.420 168.655 ;
        RECT 85.065 168.545 85.365 169.545 ;
        RECT 85.625 169.335 85.795 169.845 ;
        RECT 85.965 169.165 86.295 169.675 ;
        RECT 86.465 169.635 86.635 169.845 ;
        RECT 87.360 169.635 87.530 170.015 ;
        RECT 88.300 169.685 88.485 170.015 ;
        RECT 86.465 169.465 87.530 169.635 ;
        RECT 85.535 168.995 86.295 169.165 ;
        RECT 85.535 168.470 85.705 168.995 ;
        RECT 86.600 168.825 86.845 169.225 ;
        RECT 86.090 168.815 86.260 168.825 ;
        RECT 85.875 168.655 86.260 168.815 ;
        RECT 86.545 168.655 86.845 168.825 ;
        RECT 85.875 168.645 86.205 168.655 ;
        RECT 86.600 168.605 86.845 168.655 ;
        RECT 87.050 168.605 87.380 169.225 ;
        RECT 87.855 168.545 88.145 169.225 ;
        RECT 88.315 168.825 88.485 169.685 ;
        RECT 88.780 169.685 88.990 170.015 ;
        RECT 89.160 169.845 90.445 170.015 ;
        RECT 89.160 169.805 89.490 169.845 ;
        RECT 88.315 168.655 88.605 168.825 ;
        RECT 85.535 168.395 85.850 168.470 ;
        RECT 82.815 167.805 83.890 167.975 ;
        RECT 85.180 167.975 85.350 168.345 ;
        RECT 85.520 168.145 85.850 168.395 ;
        RECT 86.020 168.435 86.190 168.475 ;
        RECT 86.020 168.265 87.540 168.435 ;
        RECT 86.020 168.145 86.190 168.265 ;
        RECT 86.425 167.975 86.780 168.015 ;
        RECT 85.180 167.805 86.780 167.975 ;
        RECT 87.295 167.845 87.540 168.265 ;
        RECT 88.315 168.205 88.485 168.655 ;
        RECT 88.780 168.485 88.950 169.685 ;
        RECT 89.645 169.535 89.975 169.675 ;
        RECT 89.190 169.305 89.975 169.535 ;
        RECT 90.275 169.385 90.445 169.845 ;
        RECT 88.780 168.315 89.020 168.485 ;
        RECT 88.310 167.875 88.485 168.205 ;
        RECT 89.190 168.135 89.360 169.305 ;
        RECT 90.275 169.215 90.925 169.385 ;
        RECT 89.990 168.655 90.445 168.825 ;
        RECT 89.770 168.475 90.180 168.485 ;
        RECT 89.770 168.315 90.185 168.475 ;
        RECT 90.755 168.435 90.925 169.215 ;
        RECT 90.010 168.145 90.185 168.315 ;
        RECT 90.355 168.265 90.925 168.435 ;
        RECT 88.830 167.965 89.360 168.135 ;
        RECT 89.530 167.975 89.700 168.135 ;
        RECT 90.355 167.975 90.525 168.265 ;
        RECT 88.830 167.805 89.000 167.965 ;
        RECT 89.530 167.805 90.525 167.975 ;
        RECT 91.115 167.805 91.375 170.015 ;
        RECT 92.465 169.555 92.995 170.015 ;
        RECT 94.135 169.555 94.465 170.015 ;
        RECT 92.465 169.385 94.465 169.555 ;
        RECT 92.465 168.375 92.635 169.385 ;
        RECT 92.805 169.045 95.450 169.215 ;
        RECT 95.665 169.045 95.995 170.015 ;
        RECT 96.695 169.515 96.865 170.015 ;
        RECT 97.535 169.845 99.065 170.015 ;
        RECT 97.535 169.685 97.705 169.845 ;
        RECT 98.055 169.515 98.225 169.675 ;
        RECT 96.695 169.345 98.225 169.515 ;
        RECT 98.395 169.505 98.725 169.675 ;
        RECT 98.395 169.175 98.565 169.505 ;
        RECT 98.895 169.345 99.065 169.845 ;
        RECT 99.235 169.175 99.585 170.015 ;
        RECT 100.345 169.845 101.355 170.015 ;
        RECT 92.805 168.545 93.155 169.045 ;
        RECT 94.795 168.965 95.450 169.045 ;
        RECT 93.385 168.545 94.075 168.875 ;
        RECT 94.245 168.545 94.535 168.875 ;
        RECT 95.305 168.625 95.655 168.795 ;
        RECT 95.305 168.375 95.485 168.625 ;
        RECT 95.825 168.455 95.995 169.045 ;
        RECT 96.670 168.825 97.015 169.165 ;
        RECT 96.665 168.655 97.015 168.825 ;
        RECT 96.670 168.545 97.015 168.655 ;
        RECT 97.325 168.545 97.760 169.165 ;
        RECT 97.930 169.005 98.565 169.175 ;
        RECT 92.465 168.205 95.485 168.375 ;
        RECT 92.465 167.830 92.905 168.205 ;
        RECT 94.135 167.805 94.465 168.205 ;
        RECT 95.665 167.805 95.995 168.455 ;
        RECT 97.930 168.485 98.100 169.005 ;
        RECT 98.780 168.945 99.585 169.175 ;
        RECT 98.780 168.835 99.140 168.945 ;
        RECT 98.600 168.655 99.140 168.835 ;
        RECT 96.695 168.185 97.705 168.355 ;
        RECT 96.695 167.810 96.865 168.185 ;
        RECT 97.535 167.975 97.705 168.185 ;
        RECT 97.930 168.315 98.220 168.485 ;
        RECT 97.930 168.145 98.270 168.315 ;
        RECT 98.440 167.975 98.610 168.310 ;
        RECT 98.780 167.980 99.140 168.655 ;
        RECT 99.785 168.545 100.085 169.545 ;
        RECT 100.345 169.335 100.515 169.845 ;
        RECT 100.685 169.165 101.015 169.675 ;
        RECT 101.185 169.635 101.355 169.845 ;
        RECT 102.080 169.635 102.250 170.015 ;
        RECT 103.020 169.685 103.205 170.015 ;
        RECT 101.185 169.465 102.250 169.635 ;
        RECT 101.320 169.165 101.565 169.225 ;
        RECT 100.255 168.995 101.015 169.165 ;
        RECT 101.265 168.995 101.565 169.165 ;
        RECT 100.255 168.470 100.425 168.995 ;
        RECT 100.810 168.815 100.980 168.825 ;
        RECT 100.595 168.655 100.980 168.815 ;
        RECT 100.595 168.645 100.925 168.655 ;
        RECT 101.320 168.605 101.565 168.995 ;
        RECT 101.770 168.605 102.100 169.225 ;
        RECT 102.575 168.545 102.865 169.225 ;
        RECT 103.035 168.825 103.205 169.685 ;
        RECT 103.500 169.685 103.710 170.015 ;
        RECT 103.880 169.845 105.165 170.015 ;
        RECT 103.880 169.805 104.210 169.845 ;
        RECT 103.035 168.655 103.325 168.825 ;
        RECT 100.255 168.395 100.570 168.470 ;
        RECT 97.535 167.805 98.610 167.975 ;
        RECT 99.900 167.975 100.070 168.345 ;
        RECT 100.240 168.145 100.570 168.395 ;
        RECT 100.740 168.435 100.910 168.475 ;
        RECT 100.740 168.265 102.260 168.435 ;
        RECT 100.740 168.145 100.910 168.265 ;
        RECT 101.145 167.975 101.500 168.015 ;
        RECT 99.900 167.805 101.500 167.975 ;
        RECT 102.015 167.845 102.260 168.265 ;
        RECT 103.035 168.205 103.205 168.655 ;
        RECT 103.500 168.485 103.670 169.685 ;
        RECT 104.365 169.535 104.695 169.675 ;
        RECT 103.910 169.305 104.695 169.535 ;
        RECT 104.995 169.385 105.165 169.845 ;
        RECT 103.500 168.315 103.740 168.485 ;
        RECT 103.030 167.875 103.205 168.205 ;
        RECT 103.910 168.135 104.080 169.305 ;
        RECT 104.995 169.215 105.645 169.385 ;
        RECT 104.710 168.655 105.165 168.825 ;
        RECT 104.490 168.475 104.900 168.485 ;
        RECT 104.490 168.315 104.905 168.475 ;
        RECT 105.475 168.435 105.645 169.215 ;
        RECT 104.730 168.145 104.905 168.315 ;
        RECT 105.075 168.265 105.645 168.435 ;
        RECT 103.550 167.965 104.080 168.135 ;
        RECT 104.250 167.975 104.420 168.135 ;
        RECT 105.075 167.975 105.245 168.265 ;
        RECT 103.550 167.805 103.720 167.965 ;
        RECT 104.250 167.805 105.245 167.975 ;
        RECT 105.835 167.805 106.095 170.015 ;
        RECT 106.730 169.045 107.065 170.015 ;
        RECT 107.575 169.845 109.605 170.015 ;
        RECT 106.730 168.375 106.900 169.045 ;
        RECT 107.575 168.875 107.745 169.845 ;
        RECT 107.070 168.545 107.325 168.875 ;
        RECT 107.550 168.545 107.745 168.875 ;
        RECT 107.915 169.505 109.040 169.675 ;
        RECT 107.155 168.375 107.325 168.545 ;
        RECT 107.915 168.375 108.085 169.505 ;
        RECT 106.730 167.805 106.985 168.375 ;
        RECT 107.155 168.205 108.085 168.375 ;
        RECT 108.255 169.165 109.265 169.335 ;
        RECT 108.255 168.365 108.425 169.165 ;
        RECT 107.910 168.170 108.085 168.205 ;
        RECT 107.910 167.805 108.440 168.170 ;
        RECT 108.630 168.145 108.905 168.965 ;
        RECT 108.625 167.975 108.905 168.145 ;
        RECT 108.630 167.805 108.905 167.975 ;
        RECT 109.075 167.805 109.265 169.165 ;
        RECT 109.435 169.180 109.605 169.845 ;
        RECT 110.180 169.425 110.695 169.835 ;
        RECT 109.435 168.990 110.185 169.180 ;
        RECT 110.355 168.615 110.695 169.425 ;
        RECT 109.465 168.445 110.695 168.615 ;
        RECT 110.865 169.110 111.135 170.015 ;
        RECT 111.815 169.255 111.985 170.015 ;
        RECT 110.175 167.840 110.420 168.445 ;
        RECT 110.865 168.310 111.035 169.110 ;
        RECT 111.320 169.085 111.985 169.255 ;
        RECT 112.245 169.110 112.515 170.015 ;
        RECT 113.195 169.255 113.375 170.015 ;
        RECT 111.320 168.940 111.490 169.085 ;
        RECT 111.205 168.610 111.490 168.940 ;
        RECT 111.320 168.355 111.490 168.610 ;
        RECT 110.865 167.805 111.125 168.310 ;
        RECT 111.320 168.185 111.985 168.355 ;
        RECT 111.815 167.805 111.985 168.185 ;
        RECT 112.245 168.310 112.425 169.110 ;
        RECT 112.700 169.085 113.375 169.255 ;
        RECT 112.700 168.940 112.870 169.085 ;
        RECT 112.595 168.610 112.870 168.940 ;
        RECT 112.700 168.355 112.870 168.610 ;
        RECT 112.245 167.805 112.505 168.310 ;
        RECT 112.700 168.185 113.365 168.355 ;
        RECT 113.195 167.805 113.365 168.185 ;
        RECT 50.605 165.085 50.865 167.295 ;
        RECT 51.455 167.125 52.450 167.295 ;
        RECT 52.980 167.135 53.150 167.295 ;
        RECT 51.455 166.835 51.625 167.125 ;
        RECT 52.280 166.965 52.450 167.125 ;
        RECT 52.620 166.965 53.150 167.135 ;
        RECT 51.055 166.665 51.625 166.835 ;
        RECT 51.795 166.785 51.970 166.955 ;
        RECT 51.055 165.885 51.225 166.665 ;
        RECT 51.795 166.625 52.210 166.785 ;
        RECT 51.800 166.615 52.210 166.625 ;
        RECT 51.535 166.275 51.990 166.445 ;
        RECT 51.055 165.715 51.705 165.885 ;
        RECT 52.620 165.795 52.790 166.965 ;
        RECT 53.495 166.895 53.670 167.225 ;
        RECT 52.960 166.615 53.200 166.785 ;
        RECT 51.535 165.255 51.705 165.715 ;
        RECT 52.005 165.565 52.790 165.795 ;
        RECT 52.005 165.425 52.335 165.565 ;
        RECT 53.030 165.415 53.200 166.615 ;
        RECT 53.495 166.445 53.665 166.895 ;
        RECT 54.440 166.835 54.685 167.255 ;
        RECT 55.200 167.125 56.800 167.295 ;
        RECT 55.200 167.085 55.555 167.125 ;
        RECT 55.790 166.835 55.960 166.955 ;
        RECT 54.440 166.665 55.960 166.835 ;
        RECT 55.790 166.625 55.960 166.665 ;
        RECT 56.130 166.705 56.460 166.955 ;
        RECT 56.630 166.755 56.800 167.125 ;
        RECT 58.090 167.125 59.165 167.295 ;
        RECT 56.130 166.630 56.445 166.705 ;
        RECT 53.375 166.275 53.665 166.445 ;
        RECT 52.490 165.255 52.820 165.295 ;
        RECT 51.535 165.085 52.820 165.255 ;
        RECT 52.990 165.085 53.200 165.415 ;
        RECT 53.495 165.415 53.665 166.275 ;
        RECT 53.835 165.875 54.125 166.555 ;
        RECT 54.600 165.875 54.930 166.495 ;
        RECT 55.135 166.445 55.380 166.495 ;
        RECT 55.775 166.445 56.105 166.455 ;
        RECT 55.135 166.275 55.435 166.445 ;
        RECT 55.720 166.285 56.105 166.445 ;
        RECT 55.720 166.275 55.890 166.285 ;
        RECT 55.135 165.875 55.380 166.275 ;
        RECT 56.275 166.105 56.445 166.630 ;
        RECT 55.685 165.935 56.445 166.105 ;
        RECT 54.450 165.465 55.515 165.635 ;
        RECT 53.495 165.085 53.680 165.415 ;
        RECT 54.450 165.085 54.620 165.465 ;
        RECT 55.345 165.255 55.515 165.465 ;
        RECT 55.685 165.425 56.015 165.935 ;
        RECT 56.185 165.255 56.355 165.765 ;
        RECT 56.615 165.555 56.915 166.555 ;
        RECT 57.560 166.445 57.920 167.120 ;
        RECT 58.090 166.790 58.260 167.125 ;
        RECT 58.430 166.785 58.770 166.955 ;
        RECT 58.480 166.615 58.770 166.785 ;
        RECT 58.995 166.915 59.165 167.125 ;
        RECT 59.835 166.915 60.005 167.290 ;
        RECT 58.995 166.745 60.005 166.915 ;
        RECT 71.355 166.895 71.560 167.295 ;
        RECT 72.255 166.965 72.515 167.295 ;
        RECT 57.560 166.265 58.100 166.445 ;
        RECT 57.560 166.155 57.920 166.265 ;
        RECT 57.115 165.925 57.920 166.155 ;
        RECT 58.600 166.095 58.770 166.615 ;
        RECT 70.875 166.725 71.560 166.895 ;
        RECT 58.135 165.925 58.770 166.095 ;
        RECT 58.940 165.935 59.375 166.555 ;
        RECT 59.685 166.105 60.030 166.555 ;
        RECT 59.685 165.935 60.035 166.105 ;
        RECT 55.345 165.085 56.355 165.255 ;
        RECT 57.115 165.085 57.465 165.925 ;
        RECT 57.635 165.255 57.805 165.755 ;
        RECT 58.135 165.595 58.305 165.925 ;
        RECT 57.975 165.425 58.305 165.595 ;
        RECT 58.475 165.585 60.005 165.755 ;
        RECT 58.475 165.425 58.645 165.585 ;
        RECT 58.995 165.255 59.165 165.415 ;
        RECT 57.635 165.085 59.165 165.255 ;
        RECT 59.835 165.085 60.005 165.585 ;
        RECT 70.875 165.695 71.215 166.725 ;
        RECT 71.385 166.055 71.635 166.555 ;
        RECT 71.815 166.225 72.175 166.805 ;
        RECT 72.345 166.055 72.515 166.965 ;
        RECT 71.385 165.885 72.515 166.055 ;
        RECT 70.875 165.520 71.540 165.695 ;
        RECT 71.355 165.115 71.540 165.520 ;
        RECT 72.245 165.115 72.515 165.885 ;
        RECT 74.575 166.895 74.835 167.295 ;
        RECT 76.095 166.910 76.425 167.295 ;
        RECT 76.095 166.895 76.685 166.910 ;
        RECT 74.575 166.725 76.685 166.895 ;
        RECT 74.575 165.425 74.835 166.725 ;
        RECT 75.050 166.225 75.565 166.555 ;
        RECT 75.050 165.765 75.220 166.225 ;
        RECT 75.940 165.935 76.345 166.555 ;
        RECT 76.515 166.055 76.685 166.725 ;
        RECT 76.855 166.225 77.195 166.785 ;
        RECT 77.695 166.725 78.035 167.295 ;
        RECT 80.095 166.895 80.300 167.295 ;
        RECT 80.995 166.965 81.255 167.295 ;
        RECT 77.365 166.225 77.640 166.555 ;
        RECT 77.365 166.055 77.535 166.225 ;
        RECT 77.810 166.105 78.035 166.725 ;
        RECT 77.805 166.055 78.035 166.105 ;
        RECT 75.045 165.595 75.220 165.765 ;
        RECT 76.515 165.885 77.535 166.055 ;
        RECT 76.515 165.735 76.685 165.885 ;
        RECT 75.050 165.090 75.220 165.595 ;
        RECT 76.095 165.470 76.685 165.735 ;
        RECT 77.705 165.390 78.035 166.055 ;
        RECT 79.615 166.725 80.300 166.895 ;
        RECT 79.615 165.695 79.955 166.725 ;
        RECT 80.125 166.055 80.375 166.555 ;
        RECT 80.555 166.225 80.915 166.805 ;
        RECT 81.085 166.055 81.255 166.965 ;
        RECT 92.055 166.895 92.260 167.295 ;
        RECT 92.955 166.965 93.215 167.295 ;
        RECT 80.125 165.885 81.255 166.055 ;
        RECT 79.615 165.520 80.280 165.695 ;
        RECT 77.695 165.085 78.035 165.390 ;
        RECT 80.095 165.115 80.280 165.520 ;
        RECT 80.985 165.115 81.255 165.885 ;
        RECT 91.575 166.725 92.260 166.895 ;
        RECT 91.575 165.695 91.915 166.725 ;
        RECT 92.085 166.055 92.335 166.555 ;
        RECT 92.515 166.225 92.875 166.805 ;
        RECT 93.045 166.055 93.215 166.965 ;
        RECT 92.085 165.885 93.215 166.055 ;
        RECT 91.575 165.520 92.240 165.695 ;
        RECT 92.055 165.115 92.240 165.520 ;
        RECT 92.945 165.115 93.215 165.885 ;
        RECT 93.845 166.895 94.285 167.270 ;
        RECT 95.515 166.895 95.845 167.295 ;
        RECT 93.845 166.725 96.865 166.895 ;
        RECT 93.845 165.715 94.015 166.725 ;
        RECT 94.185 166.055 94.535 166.555 ;
        RECT 94.765 166.225 95.455 166.555 ;
        RECT 95.625 166.225 95.915 166.555 ;
        RECT 96.685 166.475 96.865 166.725 ;
        RECT 97.045 166.645 97.375 167.295 ;
        RECT 104.855 166.835 105.185 167.295 ;
        RECT 105.695 167.060 106.025 167.295 ;
        RECT 105.695 166.835 105.945 167.060 ;
        RECT 107.110 166.890 107.440 167.295 ;
        RECT 108.765 166.890 109.315 167.295 ;
        RECT 107.110 166.835 109.315 166.890 ;
        RECT 96.685 166.305 97.035 166.475 ;
        RECT 96.175 166.055 96.830 166.135 ;
        RECT 97.205 166.055 97.375 166.645 ;
        RECT 94.185 165.885 96.830 166.055 ;
        RECT 93.845 165.545 95.845 165.715 ;
        RECT 93.845 165.085 94.375 165.545 ;
        RECT 95.515 165.085 95.845 165.545 ;
        RECT 97.045 165.085 97.375 166.055 ;
        RECT 104.425 166.645 105.945 166.835 ;
        RECT 106.115 166.665 109.315 166.835 ;
        RECT 104.425 166.095 104.685 166.645 ;
        RECT 106.115 166.475 106.285 166.665 ;
        RECT 104.855 166.265 106.285 166.475 ;
        RECT 106.455 166.305 106.940 166.475 ;
        RECT 104.425 165.925 106.025 166.095 ;
        RECT 104.855 165.085 105.185 165.925 ;
        RECT 105.695 165.085 106.025 165.925 ;
        RECT 106.770 165.425 106.940 166.305 ;
        RECT 107.110 166.225 107.440 166.475 ;
        RECT 107.610 166.005 107.780 166.665 ;
        RECT 107.110 165.805 107.780 166.005 ;
        RECT 107.950 165.915 108.340 166.475 ;
        RECT 108.510 166.265 108.975 166.475 ;
        RECT 107.110 165.495 107.440 165.805 ;
        RECT 108.510 165.635 108.680 166.265 ;
        RECT 109.145 166.095 109.315 166.665 ;
        RECT 107.610 165.465 108.680 165.635 ;
        RECT 106.770 165.325 106.955 165.425 ;
        RECT 107.610 165.325 107.780 165.465 ;
        RECT 106.770 165.155 107.780 165.325 ;
        RECT 108.935 165.085 109.315 166.095 ;
        RECT 109.950 166.725 110.205 167.295 ;
        RECT 111.130 166.930 111.660 167.295 ;
        RECT 111.130 166.895 111.305 166.930 ;
        RECT 110.375 166.725 111.305 166.895 ;
        RECT 111.850 166.785 112.125 167.295 ;
        RECT 109.950 166.055 110.120 166.725 ;
        RECT 110.375 166.555 110.545 166.725 ;
        RECT 110.290 166.225 110.545 166.555 ;
        RECT 110.770 166.225 110.965 166.555 ;
        RECT 109.950 165.085 110.285 166.055 ;
        RECT 110.795 165.255 110.965 166.225 ;
        RECT 111.135 165.595 111.305 166.725 ;
        RECT 111.475 165.935 111.645 166.735 ;
        RECT 111.845 166.615 112.125 166.785 ;
        RECT 111.850 166.135 112.125 166.615 ;
        RECT 112.295 165.935 112.485 167.295 ;
        RECT 113.395 166.655 113.640 167.260 ;
        RECT 112.685 166.485 113.915 166.655 ;
        RECT 111.475 165.765 112.485 165.935 ;
        RECT 112.655 165.920 113.405 166.110 ;
        RECT 111.135 165.425 112.260 165.595 ;
        RECT 112.655 165.255 112.825 165.920 ;
        RECT 113.575 165.675 113.915 166.485 ;
        RECT 113.400 165.265 113.915 165.675 ;
        RECT 110.795 165.085 112.825 165.255 ;
        RECT 55.695 164.235 56.075 164.405 ;
        RECT 55.695 164.065 55.865 164.235 ;
        RECT 57.455 164.065 57.785 164.575 ;
        RECT 55.205 163.865 55.865 164.065 ;
        RECT 56.035 163.895 58.255 164.065 ;
        RECT 55.205 162.935 55.375 163.865 ;
        RECT 56.035 163.695 56.205 163.895 ;
        RECT 55.545 163.525 56.205 163.695 ;
        RECT 56.375 163.555 57.915 163.725 ;
        RECT 55.545 163.105 55.715 163.525 ;
        RECT 56.375 163.355 56.545 163.555 ;
        RECT 55.945 163.185 56.545 163.355 ;
        RECT 56.715 163.185 57.410 163.385 ;
        RECT 57.670 163.105 57.915 163.555 ;
        RECT 56.035 162.935 56.945 163.015 ;
        RECT 58.085 162.935 58.255 163.895 ;
        RECT 55.205 162.455 55.525 162.935 ;
        RECT 55.695 162.845 56.945 162.935 ;
        RECT 55.695 162.765 56.205 162.845 ;
        RECT 55.695 162.365 55.925 162.765 ;
        RECT 56.615 162.365 56.945 162.845 ;
        RECT 57.790 162.390 58.255 162.935 ;
        RECT 61.185 162.365 61.445 164.575 ;
        RECT 62.115 164.405 63.400 164.575 ;
        RECT 62.115 163.945 62.285 164.405 ;
        RECT 63.070 164.365 63.400 164.405 ;
        RECT 63.570 164.245 63.780 164.575 ;
        RECT 61.635 163.775 62.285 163.945 ;
        RECT 62.585 164.095 62.915 164.235 ;
        RECT 62.585 163.865 63.370 164.095 ;
        RECT 61.635 162.995 61.805 163.775 ;
        RECT 62.115 163.215 62.570 163.385 ;
        RECT 62.380 163.035 62.790 163.045 ;
        RECT 61.635 162.825 62.205 162.995 ;
        RECT 62.035 162.535 62.205 162.825 ;
        RECT 62.375 162.875 62.790 163.035 ;
        RECT 62.375 162.705 62.550 162.875 ;
        RECT 63.200 162.695 63.370 163.865 ;
        RECT 63.610 163.045 63.780 164.245 ;
        RECT 64.075 164.245 64.260 164.575 ;
        RECT 64.075 163.385 64.245 164.245 ;
        RECT 65.030 164.195 65.200 164.575 ;
        RECT 65.925 164.405 66.935 164.575 ;
        RECT 65.925 164.195 66.095 164.405 ;
        RECT 65.030 164.025 66.095 164.195 ;
        RECT 63.955 163.215 64.245 163.385 ;
        RECT 63.540 162.875 63.780 163.045 ;
        RECT 64.075 162.765 64.245 163.215 ;
        RECT 64.415 163.105 64.705 163.785 ;
        RECT 65.180 163.165 65.510 163.785 ;
        RECT 65.715 163.385 65.960 163.785 ;
        RECT 66.265 163.725 66.595 164.235 ;
        RECT 66.765 163.895 66.935 164.405 ;
        RECT 66.265 163.555 67.025 163.725 ;
        RECT 65.715 163.215 66.015 163.385 ;
        RECT 66.300 163.375 66.470 163.385 ;
        RECT 66.300 163.215 66.685 163.375 ;
        RECT 65.715 163.165 65.960 163.215 ;
        RECT 66.355 163.205 66.685 163.215 ;
        RECT 66.370 162.995 66.540 163.035 ;
        RECT 66.855 163.030 67.025 163.555 ;
        RECT 67.195 163.105 67.495 164.105 ;
        RECT 67.695 163.735 68.045 164.575 ;
        RECT 68.215 164.405 69.745 164.575 ;
        RECT 68.215 163.905 68.385 164.405 ;
        RECT 69.575 164.245 69.745 164.405 ;
        RECT 68.555 164.065 68.885 164.235 ;
        RECT 68.715 163.735 68.885 164.065 ;
        RECT 69.055 164.075 69.225 164.235 ;
        RECT 70.415 164.075 70.585 164.575 ;
        RECT 79.175 164.140 79.360 164.545 ;
        RECT 69.055 163.905 70.585 164.075 ;
        RECT 78.695 163.965 79.360 164.140 ;
        RECT 67.695 163.505 68.500 163.735 ;
        RECT 68.715 163.565 69.350 163.735 ;
        RECT 68.140 163.395 68.500 163.505 ;
        RECT 68.140 163.215 68.680 163.395 ;
        RECT 65.020 162.825 66.540 162.995 ;
        RECT 62.860 162.535 63.030 162.695 ;
        RECT 62.035 162.365 63.030 162.535 ;
        RECT 63.200 162.525 63.730 162.695 ;
        RECT 63.560 162.365 63.730 162.525 ;
        RECT 64.075 162.435 64.250 162.765 ;
        RECT 65.020 162.405 65.265 162.825 ;
        RECT 66.370 162.705 66.540 162.825 ;
        RECT 66.710 162.955 67.025 163.030 ;
        RECT 66.710 162.705 67.040 162.955 ;
        RECT 65.780 162.535 66.135 162.575 ;
        RECT 67.210 162.535 67.380 162.905 ;
        RECT 68.140 162.540 68.500 163.215 ;
        RECT 69.180 163.045 69.350 163.565 ;
        RECT 69.520 163.105 69.955 163.725 ;
        RECT 70.265 163.385 70.610 163.725 ;
        RECT 70.265 163.215 70.615 163.385 ;
        RECT 70.265 163.105 70.610 163.215 ;
        RECT 69.060 162.875 69.350 163.045 ;
        RECT 78.695 162.935 79.035 163.965 ;
        RECT 80.065 163.775 80.335 164.545 ;
        RECT 79.205 163.605 80.335 163.775 ;
        RECT 79.205 163.105 79.455 163.605 ;
        RECT 65.780 162.365 67.380 162.535 ;
        RECT 68.670 162.535 68.840 162.870 ;
        RECT 69.010 162.705 69.350 162.875 ;
        RECT 69.575 162.745 70.585 162.915 ;
        RECT 78.695 162.765 79.380 162.935 ;
        RECT 79.635 162.855 79.995 163.435 ;
        RECT 69.575 162.535 69.745 162.745 ;
        RECT 68.670 162.365 69.745 162.535 ;
        RECT 70.415 162.370 70.585 162.745 ;
        RECT 79.175 162.365 79.380 162.765 ;
        RECT 80.165 162.695 80.335 163.605 ;
        RECT 80.075 162.365 80.335 162.695 ;
        RECT 80.965 164.115 81.495 164.575 ;
        RECT 82.635 164.115 82.965 164.575 ;
        RECT 80.965 163.945 82.965 164.115 ;
        RECT 80.965 162.935 81.135 163.945 ;
        RECT 81.305 163.605 83.950 163.775 ;
        RECT 84.165 163.605 84.495 164.575 ;
        RECT 81.305 163.105 81.655 163.605 ;
        RECT 83.295 163.525 83.950 163.605 ;
        RECT 81.885 163.105 82.575 163.435 ;
        RECT 82.745 163.105 83.035 163.435 ;
        RECT 83.805 163.185 84.155 163.355 ;
        RECT 83.805 162.935 83.985 163.185 ;
        RECT 84.325 163.015 84.495 163.605 ;
        RECT 80.965 162.765 83.985 162.935 ;
        RECT 80.965 162.390 81.405 162.765 ;
        RECT 82.635 162.365 82.965 162.765 ;
        RECT 84.165 162.365 84.495 163.015 ;
        RECT 86.030 163.605 86.365 164.575 ;
        RECT 86.875 164.405 88.905 164.575 ;
        RECT 86.030 162.935 86.200 163.605 ;
        RECT 86.875 163.435 87.045 164.405 ;
        RECT 86.370 163.105 86.625 163.435 ;
        RECT 86.850 163.105 87.045 163.435 ;
        RECT 87.215 164.065 88.340 164.235 ;
        RECT 86.455 162.935 86.625 163.105 ;
        RECT 87.215 162.935 87.385 164.065 ;
        RECT 86.030 162.365 86.285 162.935 ;
        RECT 86.455 162.765 87.385 162.935 ;
        RECT 87.555 163.725 88.565 163.895 ;
        RECT 87.555 162.925 87.725 163.725 ;
        RECT 87.930 163.385 88.205 163.525 ;
        RECT 87.925 163.215 88.205 163.385 ;
        RECT 87.210 162.730 87.385 162.765 ;
        RECT 87.210 162.365 87.740 162.730 ;
        RECT 87.930 162.365 88.205 163.215 ;
        RECT 88.375 162.365 88.565 163.725 ;
        RECT 88.735 163.740 88.905 164.405 ;
        RECT 89.480 163.985 89.995 164.395 ;
        RECT 88.735 163.550 89.485 163.740 ;
        RECT 89.655 163.175 89.995 163.985 ;
        RECT 88.765 163.005 89.995 163.175 ;
        RECT 93.850 163.605 94.185 164.575 ;
        RECT 94.695 164.405 96.725 164.575 ;
        RECT 89.475 162.400 89.720 163.005 ;
        RECT 93.850 162.935 94.020 163.605 ;
        RECT 94.695 163.435 94.865 164.405 ;
        RECT 94.190 163.105 94.445 163.435 ;
        RECT 94.670 163.105 94.865 163.435 ;
        RECT 95.035 164.065 96.160 164.235 ;
        RECT 94.275 162.935 94.445 163.105 ;
        RECT 95.035 162.935 95.205 164.065 ;
        RECT 93.850 162.365 94.105 162.935 ;
        RECT 94.275 162.765 95.205 162.935 ;
        RECT 95.375 163.725 96.385 163.895 ;
        RECT 95.375 162.925 95.545 163.725 ;
        RECT 95.030 162.730 95.205 162.765 ;
        RECT 95.030 162.365 95.560 162.730 ;
        RECT 95.750 162.705 96.025 163.525 ;
        RECT 95.745 162.535 96.025 162.705 ;
        RECT 95.750 162.365 96.025 162.535 ;
        RECT 96.195 162.365 96.385 163.725 ;
        RECT 96.555 163.740 96.725 164.405 ;
        RECT 97.300 163.985 97.815 164.395 ;
        RECT 96.555 163.550 97.305 163.740 ;
        RECT 97.475 163.175 97.815 163.985 ;
        RECT 96.585 163.005 97.815 163.175 ;
        RECT 97.990 163.605 98.325 164.575 ;
        RECT 98.835 164.405 100.865 164.575 ;
        RECT 97.295 162.400 97.540 163.005 ;
        RECT 97.990 162.935 98.160 163.605 ;
        RECT 98.835 163.435 99.005 164.405 ;
        RECT 98.330 163.105 98.585 163.435 ;
        RECT 98.810 163.105 99.005 163.435 ;
        RECT 99.175 164.065 100.300 164.235 ;
        RECT 98.415 162.935 98.585 163.105 ;
        RECT 99.175 162.935 99.345 164.065 ;
        RECT 97.990 162.365 98.245 162.935 ;
        RECT 98.415 162.765 99.345 162.935 ;
        RECT 99.515 163.725 100.525 163.895 ;
        RECT 99.515 162.925 99.685 163.725 ;
        RECT 99.890 163.045 100.165 163.525 ;
        RECT 99.885 162.875 100.165 163.045 ;
        RECT 99.170 162.730 99.345 162.765 ;
        RECT 99.170 162.365 99.700 162.730 ;
        RECT 99.890 162.365 100.165 162.875 ;
        RECT 100.335 162.365 100.525 163.725 ;
        RECT 100.695 163.740 100.865 164.405 ;
        RECT 101.440 163.985 101.955 164.395 ;
        RECT 100.695 163.550 101.445 163.740 ;
        RECT 101.615 163.175 101.955 163.985 ;
        RECT 100.725 163.005 101.955 163.175 ;
        RECT 102.125 163.775 102.395 164.545 ;
        RECT 103.100 164.140 103.285 164.545 ;
        RECT 103.100 163.965 103.765 164.140 ;
        RECT 102.125 163.605 103.255 163.775 ;
        RECT 101.435 162.400 101.680 163.005 ;
        RECT 102.125 162.695 102.295 163.605 ;
        RECT 102.465 162.855 102.825 163.435 ;
        RECT 103.005 163.105 103.255 163.605 ;
        RECT 103.425 162.935 103.765 163.965 ;
        RECT 103.080 162.765 103.765 162.935 ;
        RECT 109.485 163.670 109.755 164.575 ;
        RECT 110.435 163.815 110.615 164.575 ;
        RECT 109.485 162.870 109.665 163.670 ;
        RECT 109.940 163.645 110.615 163.815 ;
        RECT 110.865 163.670 111.135 164.575 ;
        RECT 111.815 163.815 111.985 164.575 ;
        RECT 109.940 163.500 110.110 163.645 ;
        RECT 109.835 163.170 110.110 163.500 ;
        RECT 109.940 162.915 110.110 163.170 ;
        RECT 110.335 163.095 110.675 163.465 ;
        RECT 102.125 162.365 102.385 162.695 ;
        RECT 103.080 162.365 103.285 162.765 ;
        RECT 109.485 162.365 109.745 162.870 ;
        RECT 109.940 162.745 110.605 162.915 ;
        RECT 110.435 162.365 110.605 162.745 ;
        RECT 110.865 162.870 111.035 163.670 ;
        RECT 111.320 163.645 111.985 163.815 ;
        RECT 112.245 163.670 112.515 164.575 ;
        RECT 113.195 163.815 113.365 164.575 ;
        RECT 111.320 163.500 111.490 163.645 ;
        RECT 111.205 163.170 111.490 163.500 ;
        RECT 111.320 162.915 111.490 163.170 ;
        RECT 110.865 162.365 111.125 162.870 ;
        RECT 111.320 162.745 111.985 162.915 ;
        RECT 111.815 162.365 111.985 162.745 ;
        RECT 112.245 162.870 112.415 163.670 ;
        RECT 112.700 163.645 113.365 163.815 ;
        RECT 112.700 163.500 112.870 163.645 ;
        RECT 112.585 163.170 112.870 163.500 ;
        RECT 112.700 162.915 112.870 163.170 ;
        RECT 112.245 162.365 112.505 162.870 ;
        RECT 112.700 162.745 113.365 162.915 ;
        RECT 113.195 162.365 113.365 162.745 ;
        RECT 52.535 161.455 52.705 161.775 ;
        RECT 53.620 161.625 54.575 161.795 ;
        RECT 51.985 161.285 54.235 161.455 ;
        RECT 51.985 160.325 52.155 161.285 ;
        RECT 52.325 160.665 52.570 161.115 ;
        RECT 52.740 160.835 53.290 161.035 ;
        RECT 53.460 160.865 53.835 161.035 ;
        RECT 53.460 160.665 53.630 160.865 ;
        RECT 54.005 160.785 54.235 161.285 ;
        RECT 52.325 160.495 53.630 160.665 ;
        RECT 54.405 160.745 54.575 161.625 ;
        RECT 55.205 161.285 55.670 161.830 ;
        RECT 56.515 161.375 56.845 161.855 ;
        RECT 57.535 161.455 57.765 161.855 ;
        RECT 57.255 161.375 57.765 161.455 ;
        RECT 56.515 161.285 57.765 161.375 ;
        RECT 57.935 161.285 58.255 161.765 ;
        RECT 54.405 160.575 55.035 160.745 ;
        RECT 51.985 159.645 52.365 160.325 ;
        RECT 53.295 160.155 54.535 160.325 ;
        RECT 53.295 159.645 53.625 160.155 ;
        RECT 54.135 159.645 54.535 160.155 ;
        RECT 54.715 159.645 55.035 160.575 ;
        RECT 55.205 160.325 55.375 161.285 ;
        RECT 56.515 161.205 57.425 161.285 ;
        RECT 55.545 160.665 55.790 161.115 ;
        RECT 56.050 160.835 56.745 161.035 ;
        RECT 56.915 160.865 57.515 161.035 ;
        RECT 56.915 160.665 57.085 160.865 ;
        RECT 57.745 160.695 57.915 161.115 ;
        RECT 55.545 160.495 57.085 160.665 ;
        RECT 57.255 160.525 57.915 160.695 ;
        RECT 57.255 160.325 57.425 160.525 ;
        RECT 58.085 160.355 58.255 161.285 ;
        RECT 55.205 160.155 57.425 160.325 ;
        RECT 57.595 160.155 58.255 160.355 ;
        RECT 61.185 161.285 61.650 161.830 ;
        RECT 62.495 161.375 62.825 161.855 ;
        RECT 63.515 161.455 63.745 161.855 ;
        RECT 63.235 161.375 63.745 161.455 ;
        RECT 62.495 161.285 63.745 161.375 ;
        RECT 63.915 161.285 64.235 161.765 ;
        RECT 64.955 161.455 65.125 161.775 ;
        RECT 66.040 161.625 66.995 161.795 ;
        RECT 61.185 160.325 61.355 161.285 ;
        RECT 62.495 161.205 63.405 161.285 ;
        RECT 61.525 160.665 61.770 161.115 ;
        RECT 62.030 160.835 62.725 161.035 ;
        RECT 62.895 160.865 63.495 161.035 ;
        RECT 62.895 160.665 63.065 160.865 ;
        RECT 63.725 160.695 63.895 161.115 ;
        RECT 61.525 160.495 63.065 160.665 ;
        RECT 63.235 160.525 63.895 160.695 ;
        RECT 63.235 160.325 63.405 160.525 ;
        RECT 64.065 160.355 64.235 161.285 ;
        RECT 61.185 160.155 63.405 160.325 ;
        RECT 63.575 160.155 64.235 160.355 ;
        RECT 64.405 161.285 66.655 161.455 ;
        RECT 64.405 160.325 64.575 161.285 ;
        RECT 64.745 160.665 64.990 161.115 ;
        RECT 65.160 160.835 65.710 161.035 ;
        RECT 65.880 160.865 66.255 161.035 ;
        RECT 65.880 160.665 66.050 160.865 ;
        RECT 66.425 160.785 66.655 161.285 ;
        RECT 64.745 160.495 66.050 160.665 ;
        RECT 66.825 160.745 66.995 161.625 ;
        RECT 69.930 161.285 70.185 161.855 ;
        RECT 71.110 161.490 71.640 161.855 ;
        RECT 71.110 161.455 71.285 161.490 ;
        RECT 70.355 161.285 71.285 161.455 ;
        RECT 66.825 160.575 67.455 160.745 ;
        RECT 55.675 159.645 56.005 160.155 ;
        RECT 57.595 159.985 57.765 160.155 ;
        RECT 57.385 159.815 57.765 159.985 ;
        RECT 61.655 159.645 61.985 160.155 ;
        RECT 63.575 159.985 63.745 160.155 ;
        RECT 63.365 159.815 63.745 159.985 ;
        RECT 64.405 159.645 64.785 160.325 ;
        RECT 65.715 160.155 66.955 160.325 ;
        RECT 65.715 159.645 66.045 160.155 ;
        RECT 66.555 159.645 66.955 160.155 ;
        RECT 67.135 159.645 67.455 160.575 ;
        RECT 69.930 160.615 70.100 161.285 ;
        RECT 70.355 161.115 70.525 161.285 ;
        RECT 70.270 160.785 70.525 161.115 ;
        RECT 70.750 160.785 70.945 161.115 ;
        RECT 69.930 159.645 70.265 160.615 ;
        RECT 70.775 159.815 70.945 160.785 ;
        RECT 71.115 160.155 71.285 161.285 ;
        RECT 71.455 160.495 71.625 161.295 ;
        RECT 71.830 161.005 72.105 161.855 ;
        RECT 71.825 160.835 72.105 161.005 ;
        RECT 71.830 160.695 72.105 160.835 ;
        RECT 72.275 160.495 72.465 161.855 ;
        RECT 73.375 161.215 73.620 161.820 ;
        RECT 74.070 161.285 74.325 161.855 ;
        RECT 75.250 161.490 75.780 161.855 ;
        RECT 75.970 161.685 76.245 161.855 ;
        RECT 75.965 161.515 76.245 161.685 ;
        RECT 75.250 161.455 75.425 161.490 ;
        RECT 74.495 161.285 75.425 161.455 ;
        RECT 72.665 161.045 73.895 161.215 ;
        RECT 71.455 160.325 72.465 160.495 ;
        RECT 72.635 160.480 73.385 160.670 ;
        RECT 71.115 159.985 72.240 160.155 ;
        RECT 72.635 159.815 72.805 160.480 ;
        RECT 73.555 160.235 73.895 161.045 ;
        RECT 73.380 159.825 73.895 160.235 ;
        RECT 74.070 160.615 74.240 161.285 ;
        RECT 74.495 161.115 74.665 161.285 ;
        RECT 74.410 160.785 74.665 161.115 ;
        RECT 74.890 160.785 75.085 161.115 ;
        RECT 70.775 159.645 72.805 159.815 ;
        RECT 74.070 159.645 74.405 160.615 ;
        RECT 74.915 159.815 75.085 160.785 ;
        RECT 75.255 160.155 75.425 161.285 ;
        RECT 75.595 160.495 75.765 161.295 ;
        RECT 75.970 160.695 76.245 161.515 ;
        RECT 76.415 160.495 76.605 161.855 ;
        RECT 77.515 161.215 77.760 161.820 ;
        RECT 79.125 161.285 79.590 161.830 ;
        RECT 80.435 161.375 80.765 161.855 ;
        RECT 81.455 161.455 81.685 161.855 ;
        RECT 81.175 161.375 81.685 161.455 ;
        RECT 80.435 161.285 81.685 161.375 ;
        RECT 81.855 161.285 82.175 161.765 ;
        RECT 76.805 161.045 78.035 161.215 ;
        RECT 75.595 160.325 76.605 160.495 ;
        RECT 76.775 160.480 77.525 160.670 ;
        RECT 75.255 159.985 76.380 160.155 ;
        RECT 76.775 159.815 76.945 160.480 ;
        RECT 77.695 160.235 78.035 161.045 ;
        RECT 77.520 159.825 78.035 160.235 ;
        RECT 79.125 160.325 79.295 161.285 ;
        RECT 80.435 161.205 81.345 161.285 ;
        RECT 79.465 160.665 79.710 161.115 ;
        RECT 79.970 160.835 80.665 161.035 ;
        RECT 80.835 160.865 81.435 161.035 ;
        RECT 80.835 160.665 81.005 160.865 ;
        RECT 81.665 160.695 81.835 161.115 ;
        RECT 79.465 160.495 81.005 160.665 ;
        RECT 81.175 160.525 81.835 160.695 ;
        RECT 81.175 160.325 81.345 160.525 ;
        RECT 82.005 160.355 82.175 161.285 ;
        RECT 90.165 161.625 91.120 161.795 ;
        RECT 90.165 160.745 90.335 161.625 ;
        RECT 92.035 161.455 92.205 161.775 ;
        RECT 96.195 161.455 96.400 161.855 ;
        RECT 97.095 161.525 97.355 161.855 ;
        RECT 90.505 161.285 92.755 161.455 ;
        RECT 90.505 160.785 90.735 161.285 ;
        RECT 90.905 160.865 91.280 161.035 ;
        RECT 79.125 160.155 81.345 160.325 ;
        RECT 81.515 160.155 82.175 160.355 ;
        RECT 89.705 160.575 90.335 160.745 ;
        RECT 91.110 160.665 91.280 160.865 ;
        RECT 91.450 160.835 92.000 161.035 ;
        RECT 92.170 160.665 92.415 161.115 ;
        RECT 74.915 159.645 76.945 159.815 ;
        RECT 79.595 159.645 79.925 160.155 ;
        RECT 81.515 159.985 81.685 160.155 ;
        RECT 81.305 159.815 81.685 159.985 ;
        RECT 89.705 159.645 90.025 160.575 ;
        RECT 91.110 160.495 92.415 160.665 ;
        RECT 92.585 160.325 92.755 161.285 ;
        RECT 90.205 160.155 91.445 160.325 ;
        RECT 90.205 159.645 90.605 160.155 ;
        RECT 91.115 159.645 91.445 160.155 ;
        RECT 92.375 159.645 92.755 160.325 ;
        RECT 95.715 161.285 96.400 161.455 ;
        RECT 95.715 160.255 96.055 161.285 ;
        RECT 96.225 160.615 96.475 161.115 ;
        RECT 96.655 160.785 97.015 161.365 ;
        RECT 97.185 160.615 97.355 161.525 ;
        RECT 96.225 160.445 97.355 160.615 ;
        RECT 95.715 160.080 96.380 160.255 ;
        RECT 96.195 159.675 96.380 160.080 ;
        RECT 97.085 159.675 97.355 160.445 ;
        RECT 101.670 161.285 101.925 161.855 ;
        RECT 102.850 161.490 103.380 161.855 ;
        RECT 102.850 161.455 103.025 161.490 ;
        RECT 102.095 161.285 103.025 161.455 ;
        RECT 101.670 160.615 101.840 161.285 ;
        RECT 102.095 161.115 102.265 161.285 ;
        RECT 102.010 160.785 102.265 161.115 ;
        RECT 102.490 160.785 102.685 161.115 ;
        RECT 101.670 159.645 102.005 160.615 ;
        RECT 102.515 159.815 102.685 160.785 ;
        RECT 102.855 160.155 103.025 161.285 ;
        RECT 103.195 160.495 103.365 161.295 ;
        RECT 103.570 161.005 103.845 161.855 ;
        RECT 103.565 160.835 103.845 161.005 ;
        RECT 103.570 160.695 103.845 160.835 ;
        RECT 104.015 160.495 104.205 161.855 ;
        RECT 105.115 161.215 105.360 161.820 ;
        RECT 105.805 161.285 106.145 161.855 ;
        RECT 107.415 161.470 107.745 161.855 ;
        RECT 107.155 161.455 107.745 161.470 ;
        RECT 109.005 161.455 109.265 161.855 ;
        RECT 104.405 161.045 105.635 161.215 ;
        RECT 103.195 160.325 104.205 160.495 ;
        RECT 104.375 160.480 105.125 160.670 ;
        RECT 102.855 159.985 103.980 160.155 ;
        RECT 104.375 159.815 104.545 160.480 ;
        RECT 105.295 160.235 105.635 161.045 ;
        RECT 105.120 159.825 105.635 160.235 ;
        RECT 105.805 160.615 106.030 161.285 ;
        RECT 106.200 160.785 106.475 161.115 ;
        RECT 106.645 160.785 106.985 161.345 ;
        RECT 107.155 161.285 109.265 161.455 ;
        RECT 106.305 160.615 106.475 160.785 ;
        RECT 107.155 160.615 107.325 161.285 ;
        RECT 105.805 159.950 106.135 160.615 ;
        RECT 106.305 160.445 107.325 160.615 ;
        RECT 107.495 160.495 107.900 161.115 ;
        RECT 108.275 160.785 108.790 161.115 ;
        RECT 107.155 160.295 107.325 160.445 ;
        RECT 108.620 160.325 108.790 160.785 ;
        RECT 107.155 160.030 107.745 160.295 ;
        RECT 108.620 160.155 108.795 160.325 ;
        RECT 102.515 159.645 104.545 159.815 ;
        RECT 105.805 159.645 106.145 159.950 ;
        RECT 108.620 159.650 108.790 160.155 ;
        RECT 109.005 159.985 109.265 161.285 ;
        RECT 110.865 161.350 111.125 161.855 ;
        RECT 111.815 161.475 111.985 161.855 ;
        RECT 110.865 160.550 111.045 161.350 ;
        RECT 111.320 161.305 111.985 161.475 ;
        RECT 112.245 161.350 112.505 161.855 ;
        RECT 113.195 161.475 113.365 161.855 ;
        RECT 111.320 161.050 111.490 161.305 ;
        RECT 111.215 160.720 111.490 161.050 ;
        RECT 111.320 160.575 111.490 160.720 ;
        RECT 110.865 159.645 111.135 160.550 ;
        RECT 111.320 160.405 111.995 160.575 ;
        RECT 111.815 159.645 111.995 160.405 ;
        RECT 112.245 160.550 112.415 161.350 ;
        RECT 112.700 161.305 113.365 161.475 ;
        RECT 112.700 161.050 112.870 161.305 ;
        RECT 112.585 160.720 112.870 161.050 ;
        RECT 112.700 160.575 112.870 160.720 ;
        RECT 112.245 159.645 112.515 160.550 ;
        RECT 112.700 160.405 113.365 160.575 ;
        RECT 113.195 159.645 113.365 160.405 ;
        RECT 43.785 158.375 43.965 159.135 ;
        RECT 43.785 158.205 44.460 158.375 ;
        RECT 44.645 158.230 44.915 159.135 ;
        RECT 44.290 158.060 44.460 158.205 ;
        RECT 43.725 157.655 44.065 158.025 ;
        RECT 44.290 157.730 44.565 158.060 ;
        RECT 44.290 157.475 44.460 157.730 ;
        RECT 43.795 157.305 44.460 157.475 ;
        RECT 44.735 157.430 44.915 158.230 ;
        RECT 48.845 158.375 49.025 159.135 ;
        RECT 48.845 158.205 49.520 158.375 ;
        RECT 49.705 158.230 49.975 159.135 ;
        RECT 49.350 158.060 49.520 158.205 ;
        RECT 48.785 157.655 49.125 158.025 ;
        RECT 49.350 157.730 49.625 158.060 ;
        RECT 49.350 157.475 49.520 157.730 ;
        RECT 43.795 156.925 43.965 157.305 ;
        RECT 44.655 156.925 44.915 157.430 ;
        RECT 48.855 157.305 49.520 157.475 ;
        RECT 49.795 157.430 49.975 158.230 ;
        RECT 55.285 158.375 55.465 159.135 ;
        RECT 55.285 158.205 55.960 158.375 ;
        RECT 56.145 158.230 56.415 159.135 ;
        RECT 55.790 158.060 55.960 158.205 ;
        RECT 55.225 157.655 55.565 158.025 ;
        RECT 55.790 157.730 56.065 158.060 ;
        RECT 55.790 157.475 55.960 157.730 ;
        RECT 48.855 156.925 49.025 157.305 ;
        RECT 49.715 156.925 49.975 157.430 ;
        RECT 55.295 157.305 55.960 157.475 ;
        RECT 56.235 157.430 56.415 158.230 ;
        RECT 58.975 158.375 59.145 159.135 ;
        RECT 58.975 158.205 59.640 158.375 ;
        RECT 59.825 158.230 60.095 159.135 ;
        RECT 59.470 158.060 59.640 158.205 ;
        RECT 58.905 157.655 59.235 158.025 ;
        RECT 59.470 157.730 59.755 158.060 ;
        RECT 59.470 157.475 59.640 157.730 ;
        RECT 55.295 156.925 55.465 157.305 ;
        RECT 56.155 156.925 56.415 157.430 ;
        RECT 58.975 157.305 59.640 157.475 ;
        RECT 59.925 157.430 60.095 158.230 ;
        RECT 64.025 158.375 64.205 159.135 ;
        RECT 64.025 158.205 64.700 158.375 ;
        RECT 64.885 158.230 65.155 159.135 ;
        RECT 68.555 158.625 68.885 159.135 ;
        RECT 70.265 158.795 70.645 158.965 ;
        RECT 70.475 158.625 70.645 158.795 ;
        RECT 64.530 158.060 64.700 158.205 ;
        RECT 63.965 157.655 64.305 158.025 ;
        RECT 64.530 157.730 64.805 158.060 ;
        RECT 64.530 157.475 64.700 157.730 ;
        RECT 58.975 156.925 59.145 157.305 ;
        RECT 59.835 156.925 60.095 157.430 ;
        RECT 64.035 157.305 64.700 157.475 ;
        RECT 64.975 157.430 65.155 158.230 ;
        RECT 64.035 156.925 64.205 157.305 ;
        RECT 64.895 156.925 65.155 157.430 ;
        RECT 68.085 158.455 70.305 158.625 ;
        RECT 68.085 157.495 68.255 158.455 ;
        RECT 68.425 158.115 69.965 158.285 ;
        RECT 68.425 157.665 68.670 158.115 ;
        RECT 68.930 157.745 69.625 157.945 ;
        RECT 69.795 157.915 69.965 158.115 ;
        RECT 70.135 158.255 70.305 158.455 ;
        RECT 70.475 158.425 71.135 158.625 ;
        RECT 70.135 158.085 70.795 158.255 ;
        RECT 69.795 157.745 70.395 157.915 ;
        RECT 70.625 157.665 70.795 158.085 ;
        RECT 69.395 157.495 70.305 157.575 ;
        RECT 70.965 157.495 71.135 158.425 ;
        RECT 71.395 158.375 71.565 159.135 ;
        RECT 71.395 158.205 72.060 158.375 ;
        RECT 72.245 158.230 72.515 159.135 ;
        RECT 71.890 158.060 72.060 158.205 ;
        RECT 71.325 157.655 71.655 158.025 ;
        RECT 71.890 157.730 72.175 158.060 ;
        RECT 68.085 156.950 68.550 157.495 ;
        RECT 69.395 157.405 70.645 157.495 ;
        RECT 69.395 156.925 69.725 157.405 ;
        RECT 70.135 157.325 70.645 157.405 ;
        RECT 70.415 156.925 70.645 157.325 ;
        RECT 70.815 157.015 71.135 157.495 ;
        RECT 71.890 157.475 72.060 157.730 ;
        RECT 71.395 157.305 72.060 157.475 ;
        RECT 72.345 157.430 72.515 158.230 ;
        RECT 74.145 158.375 74.325 159.135 ;
        RECT 74.145 158.205 74.820 158.375 ;
        RECT 75.005 158.230 75.275 159.135 ;
        RECT 74.650 158.060 74.820 158.205 ;
        RECT 74.085 157.655 74.425 158.025 ;
        RECT 74.650 157.730 74.925 158.060 ;
        RECT 74.650 157.475 74.820 157.730 ;
        RECT 71.395 156.925 71.565 157.305 ;
        RECT 72.255 156.925 72.515 157.430 ;
        RECT 74.155 157.305 74.820 157.475 ;
        RECT 75.095 157.430 75.275 158.230 ;
        RECT 74.155 156.925 74.325 157.305 ;
        RECT 75.015 156.925 75.275 157.430 ;
        RECT 79.125 158.230 79.395 159.135 ;
        RECT 80.075 158.375 80.255 159.135 ;
        RECT 83.755 158.795 84.135 158.965 ;
        RECT 83.755 158.625 83.925 158.795 ;
        RECT 85.515 158.625 85.845 159.135 ;
        RECT 79.125 157.430 79.305 158.230 ;
        RECT 79.580 158.205 80.255 158.375 ;
        RECT 83.265 158.425 83.925 158.625 ;
        RECT 84.095 158.455 86.315 158.625 ;
        RECT 79.580 158.060 79.750 158.205 ;
        RECT 79.475 157.730 79.750 158.060 ;
        RECT 79.580 157.475 79.750 157.730 ;
        RECT 79.975 157.655 80.315 158.025 ;
        RECT 83.265 157.495 83.435 158.425 ;
        RECT 84.095 158.255 84.265 158.455 ;
        RECT 83.605 158.085 84.265 158.255 ;
        RECT 84.435 158.115 85.975 158.285 ;
        RECT 83.605 157.665 83.775 158.085 ;
        RECT 84.435 157.915 84.605 158.115 ;
        RECT 84.005 157.745 84.605 157.915 ;
        RECT 84.775 157.745 85.470 157.945 ;
        RECT 85.730 157.665 85.975 158.115 ;
        RECT 84.095 157.495 85.005 157.575 ;
        RECT 86.145 157.495 86.315 158.455 ;
        RECT 86.565 158.375 86.745 159.135 ;
        RECT 86.565 158.205 87.240 158.375 ;
        RECT 87.425 158.230 87.695 159.135 ;
        RECT 87.070 158.060 87.240 158.205 ;
        RECT 86.505 157.655 86.845 158.025 ;
        RECT 87.070 157.730 87.345 158.060 ;
        RECT 79.125 156.925 79.385 157.430 ;
        RECT 79.580 157.305 80.245 157.475 ;
        RECT 80.075 156.925 80.245 157.305 ;
        RECT 83.265 157.015 83.585 157.495 ;
        RECT 83.755 157.405 85.005 157.495 ;
        RECT 83.755 157.325 84.265 157.405 ;
        RECT 83.755 156.925 83.985 157.325 ;
        RECT 84.675 156.925 85.005 157.405 ;
        RECT 85.850 156.950 86.315 157.495 ;
        RECT 87.070 157.475 87.240 157.730 ;
        RECT 86.575 157.305 87.240 157.475 ;
        RECT 87.515 157.430 87.695 158.230 ;
        RECT 89.335 158.375 89.505 159.135 ;
        RECT 89.335 158.205 90.000 158.375 ;
        RECT 90.185 158.230 90.455 159.135 ;
        RECT 89.830 158.060 90.000 158.205 ;
        RECT 89.265 157.655 89.595 158.025 ;
        RECT 89.830 157.730 90.115 158.060 ;
        RECT 89.830 157.475 90.000 157.730 ;
        RECT 86.575 156.925 86.745 157.305 ;
        RECT 87.435 156.925 87.695 157.430 ;
        RECT 89.335 157.305 90.000 157.475 ;
        RECT 90.285 157.430 90.455 158.230 ;
        RECT 94.385 158.375 94.565 159.135 ;
        RECT 94.385 158.205 95.060 158.375 ;
        RECT 95.245 158.230 95.515 159.135 ;
        RECT 94.890 158.060 95.060 158.205 ;
        RECT 94.325 157.655 94.665 158.025 ;
        RECT 94.890 157.730 95.165 158.060 ;
        RECT 94.890 157.475 95.060 157.730 ;
        RECT 89.335 156.925 89.505 157.305 ;
        RECT 90.195 156.925 90.455 157.430 ;
        RECT 94.395 157.305 95.060 157.475 ;
        RECT 95.335 157.430 95.515 158.230 ;
        RECT 99.455 158.375 99.625 159.135 ;
        RECT 99.455 158.205 100.120 158.375 ;
        RECT 100.305 158.230 100.575 159.135 ;
        RECT 99.950 158.060 100.120 158.205 ;
        RECT 99.385 157.655 99.715 158.025 ;
        RECT 99.950 157.730 100.235 158.060 ;
        RECT 99.950 157.475 100.120 157.730 ;
        RECT 94.395 156.925 94.565 157.305 ;
        RECT 95.255 156.925 95.515 157.430 ;
        RECT 99.455 157.305 100.120 157.475 ;
        RECT 100.405 157.430 100.575 158.230 ;
        RECT 104.505 158.375 104.685 159.135 ;
        RECT 104.505 158.205 105.180 158.375 ;
        RECT 105.365 158.230 105.635 159.135 ;
        RECT 105.010 158.060 105.180 158.205 ;
        RECT 104.445 157.655 104.785 158.025 ;
        RECT 105.010 157.730 105.285 158.060 ;
        RECT 105.010 157.475 105.180 157.730 ;
        RECT 99.455 156.925 99.625 157.305 ;
        RECT 100.315 156.925 100.575 157.430 ;
        RECT 104.515 157.305 105.180 157.475 ;
        RECT 105.455 157.430 105.635 158.230 ;
        RECT 104.515 156.925 104.685 157.305 ;
        RECT 105.375 156.925 105.635 157.430 ;
        RECT 106.725 158.675 107.255 159.135 ;
        RECT 108.395 158.675 108.725 159.135 ;
        RECT 106.725 158.505 108.725 158.675 ;
        RECT 106.725 157.495 106.895 158.505 ;
        RECT 107.065 158.285 109.710 158.335 ;
        RECT 107.065 158.165 109.715 158.285 ;
        RECT 109.925 158.165 110.255 159.135 ;
        RECT 110.945 158.375 111.125 159.135 ;
        RECT 110.945 158.205 111.620 158.375 ;
        RECT 111.805 158.230 112.075 159.135 ;
        RECT 107.065 157.665 107.415 158.165 ;
        RECT 109.055 158.115 109.715 158.165 ;
        RECT 109.055 158.085 109.710 158.115 ;
        RECT 107.645 157.665 108.335 157.995 ;
        RECT 108.505 157.665 108.795 157.995 ;
        RECT 109.565 157.745 109.915 157.915 ;
        RECT 109.565 157.495 109.745 157.745 ;
        RECT 110.085 157.575 110.255 158.165 ;
        RECT 111.450 158.060 111.620 158.205 ;
        RECT 110.885 157.655 111.225 158.025 ;
        RECT 111.450 157.730 111.725 158.060 ;
        RECT 106.725 157.325 109.745 157.495 ;
        RECT 106.725 156.950 107.165 157.325 ;
        RECT 108.395 156.925 108.725 157.325 ;
        RECT 109.925 156.925 110.255 157.575 ;
        RECT 111.450 157.475 111.620 157.730 ;
        RECT 110.955 157.305 111.620 157.475 ;
        RECT 111.895 157.430 112.075 158.230 ;
        RECT 110.955 156.925 111.125 157.305 ;
        RECT 111.815 156.925 112.075 157.430 ;
        RECT 113.165 158.230 113.435 159.135 ;
        RECT 114.115 158.375 114.295 159.135 ;
        RECT 113.165 157.430 113.345 158.230 ;
        RECT 113.620 158.205 114.295 158.375 ;
        RECT 113.620 158.060 113.790 158.205 ;
        RECT 113.515 157.730 113.790 158.060 ;
        RECT 113.620 157.475 113.790 157.730 ;
        RECT 114.015 157.655 114.355 158.025 ;
        RECT 113.165 156.925 113.425 157.430 ;
        RECT 113.620 157.305 114.285 157.475 ;
        RECT 114.115 156.925 114.285 157.305 ;
        RECT 62.880 127.720 63.880 127.890 ;
        RECT 64.760 127.720 65.760 127.890 ;
        RECT 66.640 127.720 67.640 127.890 ;
        RECT 68.520 127.720 69.520 127.890 ;
        RECT 70.400 127.720 71.400 127.890 ;
        RECT 72.280 127.720 73.280 127.890 ;
        RECT 74.160 127.720 75.160 127.890 ;
        RECT 85.540 127.720 86.540 127.890 ;
        RECT 87.420 127.720 88.420 127.890 ;
        RECT 89.300 127.720 90.300 127.890 ;
        RECT 91.180 127.720 92.180 127.890 ;
        RECT 93.060 127.720 94.060 127.890 ;
        RECT 94.940 127.720 95.940 127.890 ;
        RECT 96.820 127.720 97.820 127.890 ;
        RECT 108.200 127.720 109.200 127.890 ;
        RECT 110.080 127.720 111.080 127.890 ;
        RECT 111.960 127.720 112.960 127.890 ;
        RECT 113.840 127.720 114.840 127.890 ;
        RECT 115.720 127.720 116.720 127.890 ;
        RECT 117.600 127.720 118.600 127.890 ;
        RECT 119.480 127.720 120.480 127.890 ;
        RECT 62.650 125.510 62.820 127.550 ;
        RECT 65.820 125.510 65.990 127.550 ;
        RECT 66.410 125.510 66.580 127.550 ;
        RECT 67.700 125.510 67.870 127.550 ;
        RECT 68.290 125.510 68.460 127.550 ;
        RECT 69.580 125.510 69.750 127.550 ;
        RECT 71.460 125.510 71.630 127.550 ;
        RECT 73.340 125.510 73.510 127.550 ;
        RECT 75.220 125.510 75.390 127.550 ;
        RECT 78.230 127.260 79.880 127.430 ;
        RECT 62.880 125.170 63.880 125.340 ;
        RECT 64.760 125.170 65.760 125.340 ;
        RECT 66.640 125.170 67.640 125.340 ;
        RECT 68.520 125.170 69.520 125.340 ;
        RECT 70.400 125.170 71.400 125.340 ;
        RECT 72.280 125.170 73.280 125.340 ;
        RECT 74.160 125.170 75.160 125.340 ;
        RECT 62.880 124.630 63.880 124.800 ;
        RECT 64.760 124.630 65.760 124.800 ;
        RECT 66.640 124.630 67.640 124.800 ;
        RECT 68.520 124.630 69.520 124.800 ;
        RECT 70.400 124.630 71.400 124.800 ;
        RECT 72.280 124.630 73.280 124.800 ;
        RECT 74.160 124.630 75.160 124.800 ;
        RECT 58.910 122.330 59.410 122.500 ;
        RECT 60.310 122.330 60.810 122.500 ;
        RECT 62.650 122.420 62.820 124.460 ;
        RECT 65.820 122.420 65.990 124.460 ;
        RECT 66.410 122.420 66.580 124.460 ;
        RECT 67.700 122.420 67.870 124.460 ;
        RECT 68.290 122.420 68.460 124.460 ;
        RECT 69.580 122.420 69.750 124.460 ;
        RECT 71.460 122.420 71.630 124.460 ;
        RECT 73.340 122.420 73.510 124.460 ;
        RECT 75.220 122.420 75.390 124.460 ;
        RECT 58.680 121.620 58.850 122.160 ;
        RECT 60.080 121.620 60.250 122.160 ;
        RECT 62.880 122.080 63.880 122.250 ;
        RECT 64.760 122.080 65.760 122.250 ;
        RECT 66.640 122.080 67.640 122.250 ;
        RECT 68.520 122.080 69.520 122.250 ;
        RECT 70.400 122.080 71.400 122.250 ;
        RECT 72.280 122.080 73.280 122.250 ;
        RECT 74.160 122.080 75.160 122.250 ;
        RECT 62.880 121.525 63.880 121.695 ;
        RECT 64.760 121.525 65.760 121.695 ;
        RECT 66.640 121.525 67.640 121.695 ;
        RECT 68.520 121.525 69.520 121.695 ;
        RECT 70.400 121.525 71.400 121.695 ;
        RECT 72.280 121.525 73.280 121.695 ;
        RECT 58.910 121.280 59.410 121.450 ;
        RECT 60.310 121.280 60.810 121.450 ;
        RECT 58.910 120.715 59.410 120.885 ;
        RECT 60.310 120.715 60.810 120.885 ;
        RECT 58.680 119.460 58.850 120.500 ;
        RECT 60.080 119.460 60.250 120.500 ;
        RECT 58.910 119.075 59.410 119.245 ;
        RECT 60.310 119.075 60.810 119.245 ;
        RECT 62.650 117.270 62.820 121.310 ;
        RECT 63.940 117.270 64.110 121.310 ;
        RECT 64.530 117.270 64.700 121.310 ;
        RECT 65.820 117.270 65.990 121.310 ;
        RECT 66.410 117.270 66.580 121.310 ;
        RECT 69.580 117.270 69.750 121.310 ;
        RECT 71.460 117.270 71.630 121.310 ;
        RECT 73.340 117.270 73.510 121.310 ;
        RECT 74.050 119.360 74.400 121.520 ;
        RECT 74.880 119.360 75.230 121.520 ;
        RECT 75.710 119.360 76.060 121.520 ;
        RECT 78.230 119.640 78.400 127.260 ;
        RECT 78.880 124.620 79.230 126.780 ;
        RECT 78.880 120.120 79.230 122.280 ;
        RECT 79.710 119.640 79.880 127.260 ;
        RECT 85.310 125.510 85.480 127.550 ;
        RECT 88.480 125.510 88.650 127.550 ;
        RECT 89.070 125.510 89.240 127.550 ;
        RECT 90.360 125.510 90.530 127.550 ;
        RECT 90.950 125.510 91.120 127.550 ;
        RECT 92.240 125.510 92.410 127.550 ;
        RECT 94.120 125.510 94.290 127.550 ;
        RECT 96.000 125.510 96.170 127.550 ;
        RECT 97.880 125.510 98.050 127.550 ;
        RECT 100.890 127.260 102.540 127.430 ;
        RECT 85.540 125.170 86.540 125.340 ;
        RECT 87.420 125.170 88.420 125.340 ;
        RECT 89.300 125.170 90.300 125.340 ;
        RECT 91.180 125.170 92.180 125.340 ;
        RECT 93.060 125.170 94.060 125.340 ;
        RECT 94.940 125.170 95.940 125.340 ;
        RECT 96.820 125.170 97.820 125.340 ;
        RECT 85.540 124.630 86.540 124.800 ;
        RECT 87.420 124.630 88.420 124.800 ;
        RECT 89.300 124.630 90.300 124.800 ;
        RECT 91.180 124.630 92.180 124.800 ;
        RECT 93.060 124.630 94.060 124.800 ;
        RECT 94.940 124.630 95.940 124.800 ;
        RECT 96.820 124.630 97.820 124.800 ;
        RECT 81.570 122.330 82.070 122.500 ;
        RECT 82.970 122.330 83.470 122.500 ;
        RECT 85.310 122.420 85.480 124.460 ;
        RECT 88.480 122.420 88.650 124.460 ;
        RECT 89.070 122.420 89.240 124.460 ;
        RECT 90.360 122.420 90.530 124.460 ;
        RECT 90.950 122.420 91.120 124.460 ;
        RECT 92.240 122.420 92.410 124.460 ;
        RECT 94.120 122.420 94.290 124.460 ;
        RECT 96.000 122.420 96.170 124.460 ;
        RECT 97.880 122.420 98.050 124.460 ;
        RECT 81.340 121.620 81.510 122.160 ;
        RECT 82.740 121.620 82.910 122.160 ;
        RECT 85.540 122.080 86.540 122.250 ;
        RECT 87.420 122.080 88.420 122.250 ;
        RECT 89.300 122.080 90.300 122.250 ;
        RECT 91.180 122.080 92.180 122.250 ;
        RECT 93.060 122.080 94.060 122.250 ;
        RECT 94.940 122.080 95.940 122.250 ;
        RECT 96.820 122.080 97.820 122.250 ;
        RECT 85.540 121.525 86.540 121.695 ;
        RECT 87.420 121.525 88.420 121.695 ;
        RECT 89.300 121.525 90.300 121.695 ;
        RECT 91.180 121.525 92.180 121.695 ;
        RECT 93.060 121.525 94.060 121.695 ;
        RECT 94.940 121.525 95.940 121.695 ;
        RECT 81.570 121.280 82.070 121.450 ;
        RECT 82.970 121.280 83.470 121.450 ;
        RECT 81.570 120.715 82.070 120.885 ;
        RECT 82.970 120.715 83.470 120.885 ;
        RECT 78.230 119.470 79.880 119.640 ;
        RECT 62.880 116.885 63.880 117.055 ;
        RECT 64.760 116.885 65.760 117.055 ;
        RECT 66.640 116.885 67.640 117.055 ;
        RECT 68.520 116.885 69.520 117.055 ;
        RECT 70.400 116.885 71.400 117.055 ;
        RECT 72.280 116.885 73.280 117.055 ;
        RECT 62.880 116.345 63.880 116.515 ;
        RECT 64.760 116.345 65.760 116.515 ;
        RECT 66.640 116.345 67.640 116.515 ;
        RECT 68.520 116.345 69.520 116.515 ;
        RECT 70.400 116.345 71.400 116.515 ;
        RECT 72.280 116.345 73.280 116.515 ;
        RECT 62.650 112.090 62.820 116.130 ;
        RECT 63.940 112.090 64.110 116.130 ;
        RECT 64.530 112.090 64.700 116.130 ;
        RECT 65.820 112.090 65.990 116.130 ;
        RECT 66.410 112.090 66.580 116.130 ;
        RECT 69.580 112.090 69.750 116.130 ;
        RECT 71.460 112.090 71.630 116.130 ;
        RECT 73.340 112.090 73.510 116.130 ;
        RECT 62.880 111.705 63.880 111.875 ;
        RECT 64.760 111.705 65.760 111.875 ;
        RECT 66.640 111.705 67.640 111.875 ;
        RECT 68.520 111.705 69.520 111.875 ;
        RECT 70.400 111.705 71.400 111.875 ;
        RECT 72.280 111.705 73.280 111.875 ;
        RECT 74.050 111.110 74.400 113.270 ;
        RECT 74.880 111.110 75.230 113.270 ;
        RECT 75.710 111.110 76.060 113.270 ;
        RECT 76.540 111.110 76.890 113.270 ;
        RECT 78.230 111.850 78.400 119.470 ;
        RECT 78.880 116.830 79.230 118.990 ;
        RECT 78.880 112.330 79.230 114.490 ;
        RECT 79.710 111.850 79.880 119.470 ;
        RECT 81.340 119.460 81.510 120.500 ;
        RECT 82.740 119.460 82.910 120.500 ;
        RECT 81.570 119.075 82.070 119.245 ;
        RECT 82.970 119.075 83.470 119.245 ;
        RECT 85.310 117.270 85.480 121.310 ;
        RECT 86.600 117.270 86.770 121.310 ;
        RECT 87.190 117.270 87.360 121.310 ;
        RECT 88.480 117.270 88.650 121.310 ;
        RECT 89.070 117.270 89.240 121.310 ;
        RECT 92.240 117.270 92.410 121.310 ;
        RECT 94.120 117.270 94.290 121.310 ;
        RECT 96.000 117.270 96.170 121.310 ;
        RECT 96.710 119.360 97.060 121.520 ;
        RECT 97.540 119.360 97.890 121.520 ;
        RECT 98.370 119.360 98.720 121.520 ;
        RECT 100.890 119.640 101.060 127.260 ;
        RECT 101.540 124.620 101.890 126.780 ;
        RECT 101.540 120.120 101.890 122.280 ;
        RECT 102.370 119.640 102.540 127.260 ;
        RECT 107.970 125.510 108.140 127.550 ;
        RECT 111.140 125.510 111.310 127.550 ;
        RECT 111.730 125.510 111.900 127.550 ;
        RECT 113.020 125.510 113.190 127.550 ;
        RECT 113.610 125.510 113.780 127.550 ;
        RECT 114.900 125.510 115.070 127.550 ;
        RECT 116.780 125.510 116.950 127.550 ;
        RECT 118.660 125.510 118.830 127.550 ;
        RECT 120.540 125.510 120.710 127.550 ;
        RECT 123.550 127.260 125.200 127.430 ;
        RECT 108.200 125.170 109.200 125.340 ;
        RECT 110.080 125.170 111.080 125.340 ;
        RECT 111.960 125.170 112.960 125.340 ;
        RECT 113.840 125.170 114.840 125.340 ;
        RECT 115.720 125.170 116.720 125.340 ;
        RECT 117.600 125.170 118.600 125.340 ;
        RECT 119.480 125.170 120.480 125.340 ;
        RECT 108.200 124.630 109.200 124.800 ;
        RECT 110.080 124.630 111.080 124.800 ;
        RECT 111.960 124.630 112.960 124.800 ;
        RECT 113.840 124.630 114.840 124.800 ;
        RECT 115.720 124.630 116.720 124.800 ;
        RECT 117.600 124.630 118.600 124.800 ;
        RECT 119.480 124.630 120.480 124.800 ;
        RECT 104.230 122.330 104.730 122.500 ;
        RECT 105.630 122.330 106.130 122.500 ;
        RECT 107.970 122.420 108.140 124.460 ;
        RECT 111.140 122.420 111.310 124.460 ;
        RECT 111.730 122.420 111.900 124.460 ;
        RECT 113.020 122.420 113.190 124.460 ;
        RECT 113.610 122.420 113.780 124.460 ;
        RECT 114.900 122.420 115.070 124.460 ;
        RECT 116.780 122.420 116.950 124.460 ;
        RECT 118.660 122.420 118.830 124.460 ;
        RECT 120.540 122.420 120.710 124.460 ;
        RECT 104.000 121.620 104.170 122.160 ;
        RECT 105.400 121.620 105.570 122.160 ;
        RECT 108.200 122.080 109.200 122.250 ;
        RECT 110.080 122.080 111.080 122.250 ;
        RECT 111.960 122.080 112.960 122.250 ;
        RECT 113.840 122.080 114.840 122.250 ;
        RECT 115.720 122.080 116.720 122.250 ;
        RECT 117.600 122.080 118.600 122.250 ;
        RECT 119.480 122.080 120.480 122.250 ;
        RECT 108.200 121.525 109.200 121.695 ;
        RECT 110.080 121.525 111.080 121.695 ;
        RECT 111.960 121.525 112.960 121.695 ;
        RECT 113.840 121.525 114.840 121.695 ;
        RECT 115.720 121.525 116.720 121.695 ;
        RECT 117.600 121.525 118.600 121.695 ;
        RECT 104.230 121.280 104.730 121.450 ;
        RECT 105.630 121.280 106.130 121.450 ;
        RECT 104.230 120.715 104.730 120.885 ;
        RECT 105.630 120.715 106.130 120.885 ;
        RECT 100.890 119.470 102.540 119.640 ;
        RECT 85.540 116.885 86.540 117.055 ;
        RECT 87.420 116.885 88.420 117.055 ;
        RECT 89.300 116.885 90.300 117.055 ;
        RECT 91.180 116.885 92.180 117.055 ;
        RECT 93.060 116.885 94.060 117.055 ;
        RECT 94.940 116.885 95.940 117.055 ;
        RECT 85.540 116.345 86.540 116.515 ;
        RECT 87.420 116.345 88.420 116.515 ;
        RECT 89.300 116.345 90.300 116.515 ;
        RECT 91.180 116.345 92.180 116.515 ;
        RECT 93.060 116.345 94.060 116.515 ;
        RECT 94.940 116.345 95.940 116.515 ;
        RECT 85.310 112.090 85.480 116.130 ;
        RECT 86.600 112.090 86.770 116.130 ;
        RECT 87.190 112.090 87.360 116.130 ;
        RECT 88.480 112.090 88.650 116.130 ;
        RECT 89.070 112.090 89.240 116.130 ;
        RECT 92.240 112.090 92.410 116.130 ;
        RECT 94.120 112.090 94.290 116.130 ;
        RECT 96.000 112.090 96.170 116.130 ;
        RECT 78.230 111.680 79.880 111.850 ;
        RECT 85.540 111.705 86.540 111.875 ;
        RECT 87.420 111.705 88.420 111.875 ;
        RECT 89.300 111.705 90.300 111.875 ;
        RECT 91.180 111.705 92.180 111.875 ;
        RECT 93.060 111.705 94.060 111.875 ;
        RECT 94.940 111.705 95.940 111.875 ;
        RECT 96.710 111.110 97.060 113.270 ;
        RECT 97.540 111.110 97.890 113.270 ;
        RECT 98.370 111.110 98.720 113.270 ;
        RECT 99.200 111.110 99.550 113.270 ;
        RECT 100.890 111.850 101.060 119.470 ;
        RECT 101.540 116.830 101.890 118.990 ;
        RECT 101.540 112.330 101.890 114.490 ;
        RECT 102.370 111.850 102.540 119.470 ;
        RECT 104.000 119.460 104.170 120.500 ;
        RECT 105.400 119.460 105.570 120.500 ;
        RECT 104.230 119.075 104.730 119.245 ;
        RECT 105.630 119.075 106.130 119.245 ;
        RECT 107.970 117.270 108.140 121.310 ;
        RECT 109.260 117.270 109.430 121.310 ;
        RECT 109.850 117.270 110.020 121.310 ;
        RECT 111.140 117.270 111.310 121.310 ;
        RECT 111.730 117.270 111.900 121.310 ;
        RECT 114.900 117.270 115.070 121.310 ;
        RECT 116.780 117.270 116.950 121.310 ;
        RECT 118.660 117.270 118.830 121.310 ;
        RECT 119.370 119.360 119.720 121.520 ;
        RECT 120.200 119.360 120.550 121.520 ;
        RECT 121.030 119.360 121.380 121.520 ;
        RECT 123.550 119.640 123.720 127.260 ;
        RECT 124.200 120.120 124.550 122.280 ;
        RECT 125.030 119.640 125.200 127.260 ;
        RECT 123.550 119.470 125.200 119.640 ;
        RECT 108.200 116.885 109.200 117.055 ;
        RECT 110.080 116.885 111.080 117.055 ;
        RECT 111.960 116.885 112.960 117.055 ;
        RECT 113.840 116.885 114.840 117.055 ;
        RECT 115.720 116.885 116.720 117.055 ;
        RECT 117.600 116.885 118.600 117.055 ;
        RECT 108.200 116.345 109.200 116.515 ;
        RECT 110.080 116.345 111.080 116.515 ;
        RECT 111.960 116.345 112.960 116.515 ;
        RECT 113.840 116.345 114.840 116.515 ;
        RECT 115.720 116.345 116.720 116.515 ;
        RECT 117.600 116.345 118.600 116.515 ;
        RECT 107.970 112.090 108.140 116.130 ;
        RECT 109.260 112.090 109.430 116.130 ;
        RECT 109.850 112.090 110.020 116.130 ;
        RECT 111.140 112.090 111.310 116.130 ;
        RECT 111.730 112.090 111.900 116.130 ;
        RECT 114.900 112.090 115.070 116.130 ;
        RECT 116.780 112.090 116.950 116.130 ;
        RECT 118.660 112.090 118.830 116.130 ;
        RECT 100.890 111.680 102.540 111.850 ;
        RECT 108.200 111.705 109.200 111.875 ;
        RECT 110.080 111.705 111.080 111.875 ;
        RECT 111.960 111.705 112.960 111.875 ;
        RECT 113.840 111.705 114.840 111.875 ;
        RECT 115.720 111.705 116.720 111.875 ;
        RECT 117.600 111.705 118.600 111.875 ;
        RECT 119.370 111.110 119.720 113.270 ;
        RECT 120.200 111.110 120.550 113.270 ;
        RECT 121.030 111.110 121.380 113.270 ;
        RECT 121.860 111.110 122.210 113.270 ;
        RECT 123.550 111.850 123.720 119.470 ;
        RECT 124.200 116.830 124.550 118.990 ;
        RECT 124.200 112.330 124.550 114.490 ;
        RECT 125.030 111.850 125.200 119.470 ;
        RECT 123.550 111.680 125.200 111.850 ;
        RECT 40.220 110.380 41.220 110.550 ;
        RECT 42.100 110.380 43.100 110.550 ;
        RECT 43.980 110.380 44.980 110.550 ;
        RECT 45.860 110.380 46.860 110.550 ;
        RECT 47.740 110.380 48.740 110.550 ;
        RECT 49.620 110.380 50.620 110.550 ;
        RECT 51.500 110.380 52.500 110.550 ;
        RECT 62.880 110.380 63.880 110.550 ;
        RECT 64.760 110.380 65.760 110.550 ;
        RECT 66.640 110.380 67.640 110.550 ;
        RECT 68.520 110.380 69.520 110.550 ;
        RECT 70.400 110.380 71.400 110.550 ;
        RECT 72.280 110.380 73.280 110.550 ;
        RECT 74.160 110.380 75.160 110.550 ;
        RECT 85.540 110.380 86.540 110.550 ;
        RECT 87.420 110.380 88.420 110.550 ;
        RECT 89.300 110.380 90.300 110.550 ;
        RECT 91.180 110.380 92.180 110.550 ;
        RECT 93.060 110.380 94.060 110.550 ;
        RECT 94.940 110.380 95.940 110.550 ;
        RECT 96.820 110.380 97.820 110.550 ;
        RECT 108.200 110.380 109.200 110.550 ;
        RECT 110.080 110.380 111.080 110.550 ;
        RECT 111.960 110.380 112.960 110.550 ;
        RECT 113.840 110.380 114.840 110.550 ;
        RECT 115.720 110.380 116.720 110.550 ;
        RECT 117.600 110.380 118.600 110.550 ;
        RECT 119.480 110.380 120.480 110.550 ;
        RECT 39.990 108.170 40.160 110.210 ;
        RECT 43.160 108.170 43.330 110.210 ;
        RECT 43.750 108.170 43.920 110.210 ;
        RECT 45.040 108.170 45.210 110.210 ;
        RECT 45.630 108.170 45.800 110.210 ;
        RECT 46.920 108.170 47.090 110.210 ;
        RECT 48.800 108.170 48.970 110.210 ;
        RECT 50.680 108.170 50.850 110.210 ;
        RECT 52.560 108.170 52.730 110.210 ;
        RECT 55.570 109.920 57.220 110.090 ;
        RECT 40.220 107.830 41.220 108.000 ;
        RECT 42.100 107.830 43.100 108.000 ;
        RECT 43.980 107.830 44.980 108.000 ;
        RECT 45.860 107.830 46.860 108.000 ;
        RECT 47.740 107.830 48.740 108.000 ;
        RECT 49.620 107.830 50.620 108.000 ;
        RECT 51.500 107.830 52.500 108.000 ;
        RECT 40.220 107.290 41.220 107.460 ;
        RECT 42.100 107.290 43.100 107.460 ;
        RECT 43.980 107.290 44.980 107.460 ;
        RECT 45.860 107.290 46.860 107.460 ;
        RECT 47.740 107.290 48.740 107.460 ;
        RECT 49.620 107.290 50.620 107.460 ;
        RECT 51.500 107.290 52.500 107.460 ;
        RECT 36.250 104.990 36.750 105.160 ;
        RECT 37.650 104.990 38.150 105.160 ;
        RECT 39.990 105.080 40.160 107.120 ;
        RECT 43.160 105.080 43.330 107.120 ;
        RECT 43.750 105.080 43.920 107.120 ;
        RECT 45.040 105.080 45.210 107.120 ;
        RECT 45.630 105.080 45.800 107.120 ;
        RECT 46.920 105.080 47.090 107.120 ;
        RECT 48.800 105.080 48.970 107.120 ;
        RECT 50.680 105.080 50.850 107.120 ;
        RECT 52.560 105.080 52.730 107.120 ;
        RECT 36.020 104.280 36.190 104.820 ;
        RECT 37.420 104.280 37.590 104.820 ;
        RECT 40.220 104.740 41.220 104.910 ;
        RECT 42.100 104.740 43.100 104.910 ;
        RECT 43.980 104.740 44.980 104.910 ;
        RECT 45.860 104.740 46.860 104.910 ;
        RECT 47.740 104.740 48.740 104.910 ;
        RECT 49.620 104.740 50.620 104.910 ;
        RECT 51.500 104.740 52.500 104.910 ;
        RECT 40.220 104.185 41.220 104.355 ;
        RECT 42.100 104.185 43.100 104.355 ;
        RECT 43.980 104.185 44.980 104.355 ;
        RECT 45.860 104.185 46.860 104.355 ;
        RECT 47.740 104.185 48.740 104.355 ;
        RECT 49.620 104.185 50.620 104.355 ;
        RECT 36.250 103.940 36.750 104.110 ;
        RECT 37.650 103.940 38.150 104.110 ;
        RECT 36.250 103.375 36.750 103.545 ;
        RECT 37.650 103.375 38.150 103.545 ;
        RECT 36.020 102.120 36.190 103.160 ;
        RECT 37.420 102.120 37.590 103.160 ;
        RECT 36.250 101.735 36.750 101.905 ;
        RECT 37.650 101.735 38.150 101.905 ;
        RECT 39.990 99.930 40.160 103.970 ;
        RECT 41.280 99.930 41.450 103.970 ;
        RECT 41.870 99.930 42.040 103.970 ;
        RECT 43.160 99.930 43.330 103.970 ;
        RECT 43.750 99.930 43.920 103.970 ;
        RECT 46.920 99.930 47.090 103.970 ;
        RECT 48.800 99.930 48.970 103.970 ;
        RECT 50.680 99.930 50.850 103.970 ;
        RECT 51.390 102.020 51.740 104.180 ;
        RECT 52.220 102.020 52.570 104.180 ;
        RECT 53.050 102.020 53.400 104.180 ;
        RECT 55.570 102.300 55.740 109.920 ;
        RECT 56.220 102.780 56.570 104.940 ;
        RECT 57.050 102.300 57.220 109.920 ;
        RECT 62.650 108.170 62.820 110.210 ;
        RECT 65.820 108.170 65.990 110.210 ;
        RECT 66.410 108.170 66.580 110.210 ;
        RECT 67.700 108.170 67.870 110.210 ;
        RECT 68.290 108.170 68.460 110.210 ;
        RECT 69.580 108.170 69.750 110.210 ;
        RECT 71.460 108.170 71.630 110.210 ;
        RECT 73.340 108.170 73.510 110.210 ;
        RECT 75.220 108.170 75.390 110.210 ;
        RECT 78.230 109.920 79.880 110.090 ;
        RECT 62.880 107.830 63.880 108.000 ;
        RECT 64.760 107.830 65.760 108.000 ;
        RECT 66.640 107.830 67.640 108.000 ;
        RECT 68.520 107.830 69.520 108.000 ;
        RECT 70.400 107.830 71.400 108.000 ;
        RECT 72.280 107.830 73.280 108.000 ;
        RECT 74.160 107.830 75.160 108.000 ;
        RECT 62.880 107.290 63.880 107.460 ;
        RECT 64.760 107.290 65.760 107.460 ;
        RECT 66.640 107.290 67.640 107.460 ;
        RECT 68.520 107.290 69.520 107.460 ;
        RECT 70.400 107.290 71.400 107.460 ;
        RECT 72.280 107.290 73.280 107.460 ;
        RECT 74.160 107.290 75.160 107.460 ;
        RECT 58.910 104.990 59.410 105.160 ;
        RECT 60.310 104.990 60.810 105.160 ;
        RECT 62.650 105.080 62.820 107.120 ;
        RECT 65.820 105.080 65.990 107.120 ;
        RECT 66.410 105.080 66.580 107.120 ;
        RECT 67.700 105.080 67.870 107.120 ;
        RECT 68.290 105.080 68.460 107.120 ;
        RECT 69.580 105.080 69.750 107.120 ;
        RECT 71.460 105.080 71.630 107.120 ;
        RECT 73.340 105.080 73.510 107.120 ;
        RECT 75.220 105.080 75.390 107.120 ;
        RECT 58.680 104.280 58.850 104.820 ;
        RECT 60.080 104.280 60.250 104.820 ;
        RECT 62.880 104.740 63.880 104.910 ;
        RECT 64.760 104.740 65.760 104.910 ;
        RECT 66.640 104.740 67.640 104.910 ;
        RECT 68.520 104.740 69.520 104.910 ;
        RECT 70.400 104.740 71.400 104.910 ;
        RECT 72.280 104.740 73.280 104.910 ;
        RECT 74.160 104.740 75.160 104.910 ;
        RECT 62.880 104.185 63.880 104.355 ;
        RECT 64.760 104.185 65.760 104.355 ;
        RECT 66.640 104.185 67.640 104.355 ;
        RECT 68.520 104.185 69.520 104.355 ;
        RECT 70.400 104.185 71.400 104.355 ;
        RECT 72.280 104.185 73.280 104.355 ;
        RECT 58.910 103.940 59.410 104.110 ;
        RECT 60.310 103.940 60.810 104.110 ;
        RECT 58.910 103.375 59.410 103.545 ;
        RECT 60.310 103.375 60.810 103.545 ;
        RECT 55.570 102.130 57.220 102.300 ;
        RECT 40.220 99.545 41.220 99.715 ;
        RECT 42.100 99.545 43.100 99.715 ;
        RECT 43.980 99.545 44.980 99.715 ;
        RECT 45.860 99.545 46.860 99.715 ;
        RECT 47.740 99.545 48.740 99.715 ;
        RECT 49.620 99.545 50.620 99.715 ;
        RECT 40.220 99.005 41.220 99.175 ;
        RECT 42.100 99.005 43.100 99.175 ;
        RECT 43.980 99.005 44.980 99.175 ;
        RECT 45.860 99.005 46.860 99.175 ;
        RECT 47.740 99.005 48.740 99.175 ;
        RECT 49.620 99.005 50.620 99.175 ;
        RECT 39.990 94.750 40.160 98.790 ;
        RECT 41.280 94.750 41.450 98.790 ;
        RECT 41.870 94.750 42.040 98.790 ;
        RECT 43.160 94.750 43.330 98.790 ;
        RECT 43.750 94.750 43.920 98.790 ;
        RECT 46.920 94.750 47.090 98.790 ;
        RECT 48.800 94.750 48.970 98.790 ;
        RECT 50.680 94.750 50.850 98.790 ;
        RECT 40.220 94.365 41.220 94.535 ;
        RECT 42.100 94.365 43.100 94.535 ;
        RECT 43.980 94.365 44.980 94.535 ;
        RECT 45.860 94.365 46.860 94.535 ;
        RECT 47.740 94.365 48.740 94.535 ;
        RECT 49.620 94.365 50.620 94.535 ;
        RECT 51.390 93.770 51.740 95.930 ;
        RECT 52.220 93.770 52.570 95.930 ;
        RECT 53.050 93.770 53.400 95.930 ;
        RECT 53.880 93.770 54.230 95.930 ;
        RECT 55.570 94.510 55.740 102.130 ;
        RECT 56.220 99.490 56.570 101.650 ;
        RECT 56.220 94.990 56.570 97.150 ;
        RECT 57.050 94.510 57.220 102.130 ;
        RECT 58.680 102.120 58.850 103.160 ;
        RECT 60.080 102.120 60.250 103.160 ;
        RECT 58.910 101.735 59.410 101.905 ;
        RECT 60.310 101.735 60.810 101.905 ;
        RECT 62.650 99.930 62.820 103.970 ;
        RECT 63.940 99.930 64.110 103.970 ;
        RECT 64.530 99.930 64.700 103.970 ;
        RECT 65.820 99.930 65.990 103.970 ;
        RECT 66.410 99.930 66.580 103.970 ;
        RECT 69.580 99.930 69.750 103.970 ;
        RECT 71.460 99.930 71.630 103.970 ;
        RECT 73.340 99.930 73.510 103.970 ;
        RECT 74.050 102.020 74.400 104.180 ;
        RECT 74.880 102.020 75.230 104.180 ;
        RECT 75.710 102.020 76.060 104.180 ;
        RECT 78.230 102.300 78.400 109.920 ;
        RECT 78.880 107.280 79.230 109.440 ;
        RECT 78.880 102.780 79.230 104.940 ;
        RECT 79.710 102.300 79.880 109.920 ;
        RECT 85.310 108.170 85.480 110.210 ;
        RECT 88.480 108.170 88.650 110.210 ;
        RECT 89.070 108.170 89.240 110.210 ;
        RECT 90.360 108.170 90.530 110.210 ;
        RECT 90.950 108.170 91.120 110.210 ;
        RECT 92.240 108.170 92.410 110.210 ;
        RECT 94.120 108.170 94.290 110.210 ;
        RECT 96.000 108.170 96.170 110.210 ;
        RECT 97.880 108.170 98.050 110.210 ;
        RECT 100.890 109.920 102.540 110.090 ;
        RECT 85.540 107.830 86.540 108.000 ;
        RECT 87.420 107.830 88.420 108.000 ;
        RECT 89.300 107.830 90.300 108.000 ;
        RECT 91.180 107.830 92.180 108.000 ;
        RECT 93.060 107.830 94.060 108.000 ;
        RECT 94.940 107.830 95.940 108.000 ;
        RECT 96.820 107.830 97.820 108.000 ;
        RECT 85.540 107.290 86.540 107.460 ;
        RECT 87.420 107.290 88.420 107.460 ;
        RECT 89.300 107.290 90.300 107.460 ;
        RECT 91.180 107.290 92.180 107.460 ;
        RECT 93.060 107.290 94.060 107.460 ;
        RECT 94.940 107.290 95.940 107.460 ;
        RECT 96.820 107.290 97.820 107.460 ;
        RECT 81.570 104.990 82.070 105.160 ;
        RECT 82.970 104.990 83.470 105.160 ;
        RECT 85.310 105.080 85.480 107.120 ;
        RECT 88.480 105.080 88.650 107.120 ;
        RECT 89.070 105.080 89.240 107.120 ;
        RECT 90.360 105.080 90.530 107.120 ;
        RECT 90.950 105.080 91.120 107.120 ;
        RECT 92.240 105.080 92.410 107.120 ;
        RECT 94.120 105.080 94.290 107.120 ;
        RECT 96.000 105.080 96.170 107.120 ;
        RECT 97.880 105.080 98.050 107.120 ;
        RECT 81.340 104.280 81.510 104.820 ;
        RECT 82.740 104.280 82.910 104.820 ;
        RECT 85.540 104.740 86.540 104.910 ;
        RECT 87.420 104.740 88.420 104.910 ;
        RECT 89.300 104.740 90.300 104.910 ;
        RECT 91.180 104.740 92.180 104.910 ;
        RECT 93.060 104.740 94.060 104.910 ;
        RECT 94.940 104.740 95.940 104.910 ;
        RECT 96.820 104.740 97.820 104.910 ;
        RECT 85.540 104.185 86.540 104.355 ;
        RECT 87.420 104.185 88.420 104.355 ;
        RECT 89.300 104.185 90.300 104.355 ;
        RECT 91.180 104.185 92.180 104.355 ;
        RECT 93.060 104.185 94.060 104.355 ;
        RECT 94.940 104.185 95.940 104.355 ;
        RECT 81.570 103.940 82.070 104.110 ;
        RECT 82.970 103.940 83.470 104.110 ;
        RECT 81.570 103.375 82.070 103.545 ;
        RECT 82.970 103.375 83.470 103.545 ;
        RECT 78.230 102.130 79.880 102.300 ;
        RECT 62.880 99.545 63.880 99.715 ;
        RECT 64.760 99.545 65.760 99.715 ;
        RECT 66.640 99.545 67.640 99.715 ;
        RECT 68.520 99.545 69.520 99.715 ;
        RECT 70.400 99.545 71.400 99.715 ;
        RECT 72.280 99.545 73.280 99.715 ;
        RECT 62.880 99.005 63.880 99.175 ;
        RECT 64.760 99.005 65.760 99.175 ;
        RECT 66.640 99.005 67.640 99.175 ;
        RECT 68.520 99.005 69.520 99.175 ;
        RECT 70.400 99.005 71.400 99.175 ;
        RECT 72.280 99.005 73.280 99.175 ;
        RECT 62.650 94.750 62.820 98.790 ;
        RECT 63.940 94.750 64.110 98.790 ;
        RECT 64.530 94.750 64.700 98.790 ;
        RECT 65.820 94.750 65.990 98.790 ;
        RECT 66.410 94.750 66.580 98.790 ;
        RECT 69.580 94.750 69.750 98.790 ;
        RECT 71.460 94.750 71.630 98.790 ;
        RECT 73.340 94.750 73.510 98.790 ;
        RECT 55.570 94.340 57.220 94.510 ;
        RECT 62.880 94.365 63.880 94.535 ;
        RECT 64.760 94.365 65.760 94.535 ;
        RECT 66.640 94.365 67.640 94.535 ;
        RECT 68.520 94.365 69.520 94.535 ;
        RECT 70.400 94.365 71.400 94.535 ;
        RECT 72.280 94.365 73.280 94.535 ;
        RECT 74.050 93.770 74.400 95.930 ;
        RECT 74.880 93.770 75.230 95.930 ;
        RECT 75.710 93.770 76.060 95.930 ;
        RECT 76.540 93.770 76.890 95.930 ;
        RECT 78.230 94.510 78.400 102.130 ;
        RECT 78.880 99.490 79.230 101.650 ;
        RECT 78.880 94.990 79.230 97.150 ;
        RECT 79.710 94.510 79.880 102.130 ;
        RECT 81.340 102.120 81.510 103.160 ;
        RECT 82.740 102.120 82.910 103.160 ;
        RECT 81.570 101.735 82.070 101.905 ;
        RECT 82.970 101.735 83.470 101.905 ;
        RECT 85.310 99.930 85.480 103.970 ;
        RECT 86.600 99.930 86.770 103.970 ;
        RECT 87.190 99.930 87.360 103.970 ;
        RECT 88.480 99.930 88.650 103.970 ;
        RECT 89.070 99.930 89.240 103.970 ;
        RECT 92.240 99.930 92.410 103.970 ;
        RECT 94.120 99.930 94.290 103.970 ;
        RECT 96.000 99.930 96.170 103.970 ;
        RECT 96.710 102.020 97.060 104.180 ;
        RECT 97.540 102.020 97.890 104.180 ;
        RECT 98.370 102.020 98.720 104.180 ;
        RECT 100.890 102.300 101.060 109.920 ;
        RECT 101.540 107.280 101.890 109.440 ;
        RECT 101.540 102.780 101.890 104.940 ;
        RECT 102.370 102.300 102.540 109.920 ;
        RECT 107.970 108.170 108.140 110.210 ;
        RECT 111.140 108.170 111.310 110.210 ;
        RECT 111.730 108.170 111.900 110.210 ;
        RECT 113.020 108.170 113.190 110.210 ;
        RECT 113.610 108.170 113.780 110.210 ;
        RECT 114.900 108.170 115.070 110.210 ;
        RECT 116.780 108.170 116.950 110.210 ;
        RECT 118.660 108.170 118.830 110.210 ;
        RECT 120.540 108.170 120.710 110.210 ;
        RECT 123.550 109.920 125.200 110.090 ;
        RECT 108.200 107.830 109.200 108.000 ;
        RECT 110.080 107.830 111.080 108.000 ;
        RECT 111.960 107.830 112.960 108.000 ;
        RECT 113.840 107.830 114.840 108.000 ;
        RECT 115.720 107.830 116.720 108.000 ;
        RECT 117.600 107.830 118.600 108.000 ;
        RECT 119.480 107.830 120.480 108.000 ;
        RECT 108.200 107.290 109.200 107.460 ;
        RECT 110.080 107.290 111.080 107.460 ;
        RECT 111.960 107.290 112.960 107.460 ;
        RECT 113.840 107.290 114.840 107.460 ;
        RECT 115.720 107.290 116.720 107.460 ;
        RECT 117.600 107.290 118.600 107.460 ;
        RECT 119.480 107.290 120.480 107.460 ;
        RECT 104.230 104.990 104.730 105.160 ;
        RECT 105.630 104.990 106.130 105.160 ;
        RECT 107.970 105.080 108.140 107.120 ;
        RECT 111.140 105.080 111.310 107.120 ;
        RECT 111.730 105.080 111.900 107.120 ;
        RECT 113.020 105.080 113.190 107.120 ;
        RECT 113.610 105.080 113.780 107.120 ;
        RECT 114.900 105.080 115.070 107.120 ;
        RECT 116.780 105.080 116.950 107.120 ;
        RECT 118.660 105.080 118.830 107.120 ;
        RECT 120.540 105.080 120.710 107.120 ;
        RECT 104.000 104.280 104.170 104.820 ;
        RECT 105.400 104.280 105.570 104.820 ;
        RECT 108.200 104.740 109.200 104.910 ;
        RECT 110.080 104.740 111.080 104.910 ;
        RECT 111.960 104.740 112.960 104.910 ;
        RECT 113.840 104.740 114.840 104.910 ;
        RECT 115.720 104.740 116.720 104.910 ;
        RECT 117.600 104.740 118.600 104.910 ;
        RECT 119.480 104.740 120.480 104.910 ;
        RECT 108.200 104.185 109.200 104.355 ;
        RECT 110.080 104.185 111.080 104.355 ;
        RECT 111.960 104.185 112.960 104.355 ;
        RECT 113.840 104.185 114.840 104.355 ;
        RECT 115.720 104.185 116.720 104.355 ;
        RECT 117.600 104.185 118.600 104.355 ;
        RECT 104.230 103.940 104.730 104.110 ;
        RECT 105.630 103.940 106.130 104.110 ;
        RECT 104.230 103.375 104.730 103.545 ;
        RECT 105.630 103.375 106.130 103.545 ;
        RECT 100.890 102.130 102.540 102.300 ;
        RECT 85.540 99.545 86.540 99.715 ;
        RECT 87.420 99.545 88.420 99.715 ;
        RECT 89.300 99.545 90.300 99.715 ;
        RECT 91.180 99.545 92.180 99.715 ;
        RECT 93.060 99.545 94.060 99.715 ;
        RECT 94.940 99.545 95.940 99.715 ;
        RECT 85.540 99.005 86.540 99.175 ;
        RECT 87.420 99.005 88.420 99.175 ;
        RECT 89.300 99.005 90.300 99.175 ;
        RECT 91.180 99.005 92.180 99.175 ;
        RECT 93.060 99.005 94.060 99.175 ;
        RECT 94.940 99.005 95.940 99.175 ;
        RECT 85.310 94.750 85.480 98.790 ;
        RECT 86.600 94.750 86.770 98.790 ;
        RECT 87.190 94.750 87.360 98.790 ;
        RECT 88.480 94.750 88.650 98.790 ;
        RECT 89.070 94.750 89.240 98.790 ;
        RECT 92.240 94.750 92.410 98.790 ;
        RECT 94.120 94.750 94.290 98.790 ;
        RECT 96.000 94.750 96.170 98.790 ;
        RECT 78.230 94.340 79.880 94.510 ;
        RECT 85.540 94.365 86.540 94.535 ;
        RECT 87.420 94.365 88.420 94.535 ;
        RECT 89.300 94.365 90.300 94.535 ;
        RECT 91.180 94.365 92.180 94.535 ;
        RECT 93.060 94.365 94.060 94.535 ;
        RECT 94.940 94.365 95.940 94.535 ;
        RECT 96.710 93.770 97.060 95.930 ;
        RECT 97.540 93.770 97.890 95.930 ;
        RECT 98.370 93.770 98.720 95.930 ;
        RECT 99.200 93.770 99.550 95.930 ;
        RECT 100.890 94.510 101.060 102.130 ;
        RECT 101.540 99.490 101.890 101.650 ;
        RECT 101.540 94.990 101.890 97.150 ;
        RECT 102.370 94.510 102.540 102.130 ;
        RECT 104.000 102.120 104.170 103.160 ;
        RECT 105.400 102.120 105.570 103.160 ;
        RECT 104.230 101.735 104.730 101.905 ;
        RECT 105.630 101.735 106.130 101.905 ;
        RECT 107.970 99.930 108.140 103.970 ;
        RECT 109.260 99.930 109.430 103.970 ;
        RECT 109.850 99.930 110.020 103.970 ;
        RECT 111.140 99.930 111.310 103.970 ;
        RECT 111.730 99.930 111.900 103.970 ;
        RECT 114.900 99.930 115.070 103.970 ;
        RECT 116.780 99.930 116.950 103.970 ;
        RECT 118.660 99.930 118.830 103.970 ;
        RECT 119.370 102.020 119.720 104.180 ;
        RECT 120.200 102.020 120.550 104.180 ;
        RECT 121.030 102.020 121.380 104.180 ;
        RECT 123.550 102.300 123.720 109.920 ;
        RECT 124.200 107.280 124.550 109.440 ;
        RECT 124.200 102.780 124.550 104.940 ;
        RECT 125.030 102.300 125.200 109.920 ;
        RECT 123.550 102.130 125.200 102.300 ;
        RECT 108.200 99.545 109.200 99.715 ;
        RECT 110.080 99.545 111.080 99.715 ;
        RECT 111.960 99.545 112.960 99.715 ;
        RECT 113.840 99.545 114.840 99.715 ;
        RECT 115.720 99.545 116.720 99.715 ;
        RECT 117.600 99.545 118.600 99.715 ;
        RECT 108.200 99.005 109.200 99.175 ;
        RECT 110.080 99.005 111.080 99.175 ;
        RECT 111.960 99.005 112.960 99.175 ;
        RECT 113.840 99.005 114.840 99.175 ;
        RECT 115.720 99.005 116.720 99.175 ;
        RECT 117.600 99.005 118.600 99.175 ;
        RECT 107.970 94.750 108.140 98.790 ;
        RECT 109.260 94.750 109.430 98.790 ;
        RECT 109.850 94.750 110.020 98.790 ;
        RECT 111.140 94.750 111.310 98.790 ;
        RECT 111.730 94.750 111.900 98.790 ;
        RECT 114.900 94.750 115.070 98.790 ;
        RECT 116.780 94.750 116.950 98.790 ;
        RECT 118.660 94.750 118.830 98.790 ;
        RECT 100.890 94.340 102.540 94.510 ;
        RECT 108.200 94.365 109.200 94.535 ;
        RECT 110.080 94.365 111.080 94.535 ;
        RECT 111.960 94.365 112.960 94.535 ;
        RECT 113.840 94.365 114.840 94.535 ;
        RECT 115.720 94.365 116.720 94.535 ;
        RECT 117.600 94.365 118.600 94.535 ;
        RECT 119.370 93.770 119.720 95.930 ;
        RECT 120.200 93.770 120.550 95.930 ;
        RECT 121.030 93.770 121.380 95.930 ;
        RECT 121.860 93.770 122.210 95.930 ;
        RECT 123.550 94.510 123.720 102.130 ;
        RECT 124.200 99.490 124.550 101.650 ;
        RECT 124.200 94.990 124.550 97.150 ;
        RECT 125.030 94.510 125.200 102.130 ;
        RECT 123.550 94.340 125.200 94.510 ;
        RECT 40.220 93.040 41.220 93.210 ;
        RECT 42.100 93.040 43.100 93.210 ;
        RECT 43.980 93.040 44.980 93.210 ;
        RECT 45.860 93.040 46.860 93.210 ;
        RECT 47.740 93.040 48.740 93.210 ;
        RECT 49.620 93.040 50.620 93.210 ;
        RECT 51.500 93.040 52.500 93.210 ;
        RECT 62.880 93.040 63.880 93.210 ;
        RECT 64.760 93.040 65.760 93.210 ;
        RECT 66.640 93.040 67.640 93.210 ;
        RECT 68.520 93.040 69.520 93.210 ;
        RECT 70.400 93.040 71.400 93.210 ;
        RECT 72.280 93.040 73.280 93.210 ;
        RECT 74.160 93.040 75.160 93.210 ;
        RECT 85.540 93.040 86.540 93.210 ;
        RECT 87.420 93.040 88.420 93.210 ;
        RECT 89.300 93.040 90.300 93.210 ;
        RECT 91.180 93.040 92.180 93.210 ;
        RECT 93.060 93.040 94.060 93.210 ;
        RECT 94.940 93.040 95.940 93.210 ;
        RECT 96.820 93.040 97.820 93.210 ;
        RECT 108.200 93.040 109.200 93.210 ;
        RECT 110.080 93.040 111.080 93.210 ;
        RECT 111.960 93.040 112.960 93.210 ;
        RECT 113.840 93.040 114.840 93.210 ;
        RECT 115.720 93.040 116.720 93.210 ;
        RECT 117.600 93.040 118.600 93.210 ;
        RECT 119.480 93.040 120.480 93.210 ;
        RECT 39.990 90.830 40.160 92.870 ;
        RECT 43.160 90.830 43.330 92.870 ;
        RECT 43.750 90.830 43.920 92.870 ;
        RECT 45.040 90.830 45.210 92.870 ;
        RECT 45.630 90.830 45.800 92.870 ;
        RECT 46.920 90.830 47.090 92.870 ;
        RECT 48.800 90.830 48.970 92.870 ;
        RECT 50.680 90.830 50.850 92.870 ;
        RECT 52.560 90.830 52.730 92.870 ;
        RECT 55.570 92.580 57.220 92.750 ;
        RECT 40.220 90.490 41.220 90.660 ;
        RECT 42.100 90.490 43.100 90.660 ;
        RECT 43.980 90.490 44.980 90.660 ;
        RECT 45.860 90.490 46.860 90.660 ;
        RECT 47.740 90.490 48.740 90.660 ;
        RECT 49.620 90.490 50.620 90.660 ;
        RECT 51.500 90.490 52.500 90.660 ;
        RECT 40.220 89.950 41.220 90.120 ;
        RECT 42.100 89.950 43.100 90.120 ;
        RECT 43.980 89.950 44.980 90.120 ;
        RECT 45.860 89.950 46.860 90.120 ;
        RECT 47.740 89.950 48.740 90.120 ;
        RECT 49.620 89.950 50.620 90.120 ;
        RECT 51.500 89.950 52.500 90.120 ;
        RECT 36.250 87.650 36.750 87.820 ;
        RECT 37.650 87.650 38.150 87.820 ;
        RECT 39.990 87.740 40.160 89.780 ;
        RECT 43.160 87.740 43.330 89.780 ;
        RECT 43.750 87.740 43.920 89.780 ;
        RECT 45.040 87.740 45.210 89.780 ;
        RECT 45.630 87.740 45.800 89.780 ;
        RECT 46.920 87.740 47.090 89.780 ;
        RECT 48.800 87.740 48.970 89.780 ;
        RECT 50.680 87.740 50.850 89.780 ;
        RECT 52.560 87.740 52.730 89.780 ;
        RECT 36.020 86.940 36.190 87.480 ;
        RECT 37.420 86.940 37.590 87.480 ;
        RECT 40.220 87.400 41.220 87.570 ;
        RECT 42.100 87.400 43.100 87.570 ;
        RECT 43.980 87.400 44.980 87.570 ;
        RECT 45.860 87.400 46.860 87.570 ;
        RECT 47.740 87.400 48.740 87.570 ;
        RECT 49.620 87.400 50.620 87.570 ;
        RECT 51.500 87.400 52.500 87.570 ;
        RECT 40.220 86.845 41.220 87.015 ;
        RECT 42.100 86.845 43.100 87.015 ;
        RECT 43.980 86.845 44.980 87.015 ;
        RECT 45.860 86.845 46.860 87.015 ;
        RECT 47.740 86.845 48.740 87.015 ;
        RECT 49.620 86.845 50.620 87.015 ;
        RECT 36.250 86.600 36.750 86.770 ;
        RECT 37.650 86.600 38.150 86.770 ;
        RECT 36.250 86.035 36.750 86.205 ;
        RECT 37.650 86.035 38.150 86.205 ;
        RECT 36.020 84.780 36.190 85.820 ;
        RECT 37.420 84.780 37.590 85.820 ;
        RECT 36.250 84.395 36.750 84.565 ;
        RECT 37.650 84.395 38.150 84.565 ;
        RECT 39.990 82.590 40.160 86.630 ;
        RECT 41.280 82.590 41.450 86.630 ;
        RECT 41.870 82.590 42.040 86.630 ;
        RECT 43.160 82.590 43.330 86.630 ;
        RECT 43.750 82.590 43.920 86.630 ;
        RECT 46.920 82.590 47.090 86.630 ;
        RECT 48.800 82.590 48.970 86.630 ;
        RECT 50.680 82.590 50.850 86.630 ;
        RECT 51.390 84.680 51.740 86.840 ;
        RECT 52.220 84.680 52.570 86.840 ;
        RECT 53.050 84.680 53.400 86.840 ;
        RECT 55.570 84.960 55.740 92.580 ;
        RECT 56.220 89.940 56.570 92.100 ;
        RECT 56.220 85.440 56.570 87.600 ;
        RECT 57.050 84.960 57.220 92.580 ;
        RECT 62.650 90.830 62.820 92.870 ;
        RECT 65.820 90.830 65.990 92.870 ;
        RECT 66.410 90.830 66.580 92.870 ;
        RECT 67.700 90.830 67.870 92.870 ;
        RECT 68.290 90.830 68.460 92.870 ;
        RECT 69.580 90.830 69.750 92.870 ;
        RECT 71.460 90.830 71.630 92.870 ;
        RECT 73.340 90.830 73.510 92.870 ;
        RECT 75.220 90.830 75.390 92.870 ;
        RECT 78.230 92.580 79.880 92.750 ;
        RECT 62.880 90.490 63.880 90.660 ;
        RECT 64.760 90.490 65.760 90.660 ;
        RECT 66.640 90.490 67.640 90.660 ;
        RECT 68.520 90.490 69.520 90.660 ;
        RECT 70.400 90.490 71.400 90.660 ;
        RECT 72.280 90.490 73.280 90.660 ;
        RECT 74.160 90.490 75.160 90.660 ;
        RECT 62.880 89.950 63.880 90.120 ;
        RECT 64.760 89.950 65.760 90.120 ;
        RECT 66.640 89.950 67.640 90.120 ;
        RECT 68.520 89.950 69.520 90.120 ;
        RECT 70.400 89.950 71.400 90.120 ;
        RECT 72.280 89.950 73.280 90.120 ;
        RECT 74.160 89.950 75.160 90.120 ;
        RECT 58.910 87.650 59.410 87.820 ;
        RECT 60.310 87.650 60.810 87.820 ;
        RECT 62.650 87.740 62.820 89.780 ;
        RECT 65.820 87.740 65.990 89.780 ;
        RECT 66.410 87.740 66.580 89.780 ;
        RECT 67.700 87.740 67.870 89.780 ;
        RECT 68.290 87.740 68.460 89.780 ;
        RECT 69.580 87.740 69.750 89.780 ;
        RECT 71.460 87.740 71.630 89.780 ;
        RECT 73.340 87.740 73.510 89.780 ;
        RECT 75.220 87.740 75.390 89.780 ;
        RECT 58.680 86.940 58.850 87.480 ;
        RECT 60.080 86.940 60.250 87.480 ;
        RECT 62.880 87.400 63.880 87.570 ;
        RECT 64.760 87.400 65.760 87.570 ;
        RECT 66.640 87.400 67.640 87.570 ;
        RECT 68.520 87.400 69.520 87.570 ;
        RECT 70.400 87.400 71.400 87.570 ;
        RECT 72.280 87.400 73.280 87.570 ;
        RECT 74.160 87.400 75.160 87.570 ;
        RECT 62.880 86.845 63.880 87.015 ;
        RECT 64.760 86.845 65.760 87.015 ;
        RECT 66.640 86.845 67.640 87.015 ;
        RECT 68.520 86.845 69.520 87.015 ;
        RECT 70.400 86.845 71.400 87.015 ;
        RECT 72.280 86.845 73.280 87.015 ;
        RECT 58.910 86.600 59.410 86.770 ;
        RECT 60.310 86.600 60.810 86.770 ;
        RECT 58.910 86.035 59.410 86.205 ;
        RECT 60.310 86.035 60.810 86.205 ;
        RECT 55.570 84.790 57.220 84.960 ;
        RECT 40.220 82.205 41.220 82.375 ;
        RECT 42.100 82.205 43.100 82.375 ;
        RECT 43.980 82.205 44.980 82.375 ;
        RECT 45.860 82.205 46.860 82.375 ;
        RECT 47.740 82.205 48.740 82.375 ;
        RECT 49.620 82.205 50.620 82.375 ;
        RECT 40.220 81.665 41.220 81.835 ;
        RECT 42.100 81.665 43.100 81.835 ;
        RECT 43.980 81.665 44.980 81.835 ;
        RECT 45.860 81.665 46.860 81.835 ;
        RECT 47.740 81.665 48.740 81.835 ;
        RECT 49.620 81.665 50.620 81.835 ;
        RECT 39.990 77.410 40.160 81.450 ;
        RECT 41.280 77.410 41.450 81.450 ;
        RECT 41.870 77.410 42.040 81.450 ;
        RECT 43.160 77.410 43.330 81.450 ;
        RECT 43.750 77.410 43.920 81.450 ;
        RECT 46.920 77.410 47.090 81.450 ;
        RECT 48.800 77.410 48.970 81.450 ;
        RECT 50.680 77.410 50.850 81.450 ;
        RECT 40.220 77.025 41.220 77.195 ;
        RECT 42.100 77.025 43.100 77.195 ;
        RECT 43.980 77.025 44.980 77.195 ;
        RECT 45.860 77.025 46.860 77.195 ;
        RECT 47.740 77.025 48.740 77.195 ;
        RECT 49.620 77.025 50.620 77.195 ;
        RECT 51.390 76.430 51.740 78.590 ;
        RECT 52.220 76.430 52.570 78.590 ;
        RECT 53.050 76.430 53.400 78.590 ;
        RECT 53.880 76.430 54.230 78.590 ;
        RECT 55.570 77.170 55.740 84.790 ;
        RECT 56.220 82.150 56.570 84.310 ;
        RECT 56.220 77.650 56.570 79.810 ;
        RECT 57.050 77.170 57.220 84.790 ;
        RECT 58.680 84.780 58.850 85.820 ;
        RECT 60.080 84.780 60.250 85.820 ;
        RECT 58.910 84.395 59.410 84.565 ;
        RECT 60.310 84.395 60.810 84.565 ;
        RECT 62.650 82.590 62.820 86.630 ;
        RECT 63.940 82.590 64.110 86.630 ;
        RECT 64.530 82.590 64.700 86.630 ;
        RECT 65.820 82.590 65.990 86.630 ;
        RECT 66.410 82.590 66.580 86.630 ;
        RECT 69.580 82.590 69.750 86.630 ;
        RECT 71.460 82.590 71.630 86.630 ;
        RECT 73.340 82.590 73.510 86.630 ;
        RECT 74.050 84.680 74.400 86.840 ;
        RECT 74.880 84.680 75.230 86.840 ;
        RECT 75.710 84.680 76.060 86.840 ;
        RECT 78.230 84.960 78.400 92.580 ;
        RECT 78.880 89.940 79.230 92.100 ;
        RECT 78.880 85.440 79.230 87.600 ;
        RECT 79.710 84.960 79.880 92.580 ;
        RECT 85.310 90.830 85.480 92.870 ;
        RECT 88.480 90.830 88.650 92.870 ;
        RECT 89.070 90.830 89.240 92.870 ;
        RECT 90.360 90.830 90.530 92.870 ;
        RECT 90.950 90.830 91.120 92.870 ;
        RECT 92.240 90.830 92.410 92.870 ;
        RECT 94.120 90.830 94.290 92.870 ;
        RECT 96.000 90.830 96.170 92.870 ;
        RECT 97.880 90.830 98.050 92.870 ;
        RECT 100.890 92.580 102.540 92.750 ;
        RECT 85.540 90.490 86.540 90.660 ;
        RECT 87.420 90.490 88.420 90.660 ;
        RECT 89.300 90.490 90.300 90.660 ;
        RECT 91.180 90.490 92.180 90.660 ;
        RECT 93.060 90.490 94.060 90.660 ;
        RECT 94.940 90.490 95.940 90.660 ;
        RECT 96.820 90.490 97.820 90.660 ;
        RECT 85.540 89.950 86.540 90.120 ;
        RECT 87.420 89.950 88.420 90.120 ;
        RECT 89.300 89.950 90.300 90.120 ;
        RECT 91.180 89.950 92.180 90.120 ;
        RECT 93.060 89.950 94.060 90.120 ;
        RECT 94.940 89.950 95.940 90.120 ;
        RECT 96.820 89.950 97.820 90.120 ;
        RECT 81.570 87.650 82.070 87.820 ;
        RECT 82.970 87.650 83.470 87.820 ;
        RECT 85.310 87.740 85.480 89.780 ;
        RECT 88.480 87.740 88.650 89.780 ;
        RECT 89.070 87.740 89.240 89.780 ;
        RECT 90.360 87.740 90.530 89.780 ;
        RECT 90.950 87.740 91.120 89.780 ;
        RECT 92.240 87.740 92.410 89.780 ;
        RECT 94.120 87.740 94.290 89.780 ;
        RECT 96.000 87.740 96.170 89.780 ;
        RECT 97.880 87.740 98.050 89.780 ;
        RECT 81.340 86.940 81.510 87.480 ;
        RECT 82.740 86.940 82.910 87.480 ;
        RECT 85.540 87.400 86.540 87.570 ;
        RECT 87.420 87.400 88.420 87.570 ;
        RECT 89.300 87.400 90.300 87.570 ;
        RECT 91.180 87.400 92.180 87.570 ;
        RECT 93.060 87.400 94.060 87.570 ;
        RECT 94.940 87.400 95.940 87.570 ;
        RECT 96.820 87.400 97.820 87.570 ;
        RECT 85.540 86.845 86.540 87.015 ;
        RECT 87.420 86.845 88.420 87.015 ;
        RECT 89.300 86.845 90.300 87.015 ;
        RECT 91.180 86.845 92.180 87.015 ;
        RECT 93.060 86.845 94.060 87.015 ;
        RECT 94.940 86.845 95.940 87.015 ;
        RECT 81.570 86.600 82.070 86.770 ;
        RECT 82.970 86.600 83.470 86.770 ;
        RECT 81.570 86.035 82.070 86.205 ;
        RECT 82.970 86.035 83.470 86.205 ;
        RECT 78.230 84.790 79.880 84.960 ;
        RECT 62.880 82.205 63.880 82.375 ;
        RECT 64.760 82.205 65.760 82.375 ;
        RECT 66.640 82.205 67.640 82.375 ;
        RECT 68.520 82.205 69.520 82.375 ;
        RECT 70.400 82.205 71.400 82.375 ;
        RECT 72.280 82.205 73.280 82.375 ;
        RECT 62.880 81.665 63.880 81.835 ;
        RECT 64.760 81.665 65.760 81.835 ;
        RECT 66.640 81.665 67.640 81.835 ;
        RECT 68.520 81.665 69.520 81.835 ;
        RECT 70.400 81.665 71.400 81.835 ;
        RECT 72.280 81.665 73.280 81.835 ;
        RECT 62.650 77.410 62.820 81.450 ;
        RECT 63.940 77.410 64.110 81.450 ;
        RECT 64.530 77.410 64.700 81.450 ;
        RECT 65.820 77.410 65.990 81.450 ;
        RECT 66.410 77.410 66.580 81.450 ;
        RECT 69.580 77.410 69.750 81.450 ;
        RECT 71.460 77.410 71.630 81.450 ;
        RECT 73.340 77.410 73.510 81.450 ;
        RECT 55.570 77.000 57.220 77.170 ;
        RECT 62.880 77.025 63.880 77.195 ;
        RECT 64.760 77.025 65.760 77.195 ;
        RECT 66.640 77.025 67.640 77.195 ;
        RECT 68.520 77.025 69.520 77.195 ;
        RECT 70.400 77.025 71.400 77.195 ;
        RECT 72.280 77.025 73.280 77.195 ;
        RECT 74.050 76.430 74.400 78.590 ;
        RECT 74.880 76.430 75.230 78.590 ;
        RECT 75.710 76.430 76.060 78.590 ;
        RECT 76.540 76.430 76.890 78.590 ;
        RECT 78.230 77.170 78.400 84.790 ;
        RECT 78.880 82.150 79.230 84.310 ;
        RECT 78.880 77.650 79.230 79.810 ;
        RECT 79.710 77.170 79.880 84.790 ;
        RECT 81.340 84.780 81.510 85.820 ;
        RECT 82.740 84.780 82.910 85.820 ;
        RECT 81.570 84.395 82.070 84.565 ;
        RECT 82.970 84.395 83.470 84.565 ;
        RECT 85.310 82.590 85.480 86.630 ;
        RECT 86.600 82.590 86.770 86.630 ;
        RECT 87.190 82.590 87.360 86.630 ;
        RECT 88.480 82.590 88.650 86.630 ;
        RECT 89.070 82.590 89.240 86.630 ;
        RECT 92.240 82.590 92.410 86.630 ;
        RECT 94.120 82.590 94.290 86.630 ;
        RECT 96.000 82.590 96.170 86.630 ;
        RECT 96.710 84.680 97.060 86.840 ;
        RECT 97.540 84.680 97.890 86.840 ;
        RECT 98.370 84.680 98.720 86.840 ;
        RECT 100.890 84.960 101.060 92.580 ;
        RECT 101.540 89.940 101.890 92.100 ;
        RECT 101.540 85.440 101.890 87.600 ;
        RECT 102.370 84.960 102.540 92.580 ;
        RECT 107.970 90.830 108.140 92.870 ;
        RECT 111.140 90.830 111.310 92.870 ;
        RECT 111.730 90.830 111.900 92.870 ;
        RECT 113.020 90.830 113.190 92.870 ;
        RECT 113.610 90.830 113.780 92.870 ;
        RECT 114.900 90.830 115.070 92.870 ;
        RECT 116.780 90.830 116.950 92.870 ;
        RECT 118.660 90.830 118.830 92.870 ;
        RECT 120.540 90.830 120.710 92.870 ;
        RECT 123.550 92.580 125.200 92.750 ;
        RECT 108.200 90.490 109.200 90.660 ;
        RECT 110.080 90.490 111.080 90.660 ;
        RECT 111.960 90.490 112.960 90.660 ;
        RECT 113.840 90.490 114.840 90.660 ;
        RECT 115.720 90.490 116.720 90.660 ;
        RECT 117.600 90.490 118.600 90.660 ;
        RECT 119.480 90.490 120.480 90.660 ;
        RECT 108.200 89.950 109.200 90.120 ;
        RECT 110.080 89.950 111.080 90.120 ;
        RECT 111.960 89.950 112.960 90.120 ;
        RECT 113.840 89.950 114.840 90.120 ;
        RECT 115.720 89.950 116.720 90.120 ;
        RECT 117.600 89.950 118.600 90.120 ;
        RECT 119.480 89.950 120.480 90.120 ;
        RECT 104.230 87.650 104.730 87.820 ;
        RECT 105.630 87.650 106.130 87.820 ;
        RECT 107.970 87.740 108.140 89.780 ;
        RECT 111.140 87.740 111.310 89.780 ;
        RECT 111.730 87.740 111.900 89.780 ;
        RECT 113.020 87.740 113.190 89.780 ;
        RECT 113.610 87.740 113.780 89.780 ;
        RECT 114.900 87.740 115.070 89.780 ;
        RECT 116.780 87.740 116.950 89.780 ;
        RECT 118.660 87.740 118.830 89.780 ;
        RECT 120.540 87.740 120.710 89.780 ;
        RECT 104.000 86.940 104.170 87.480 ;
        RECT 105.400 86.940 105.570 87.480 ;
        RECT 108.200 87.400 109.200 87.570 ;
        RECT 110.080 87.400 111.080 87.570 ;
        RECT 111.960 87.400 112.960 87.570 ;
        RECT 113.840 87.400 114.840 87.570 ;
        RECT 115.720 87.400 116.720 87.570 ;
        RECT 117.600 87.400 118.600 87.570 ;
        RECT 119.480 87.400 120.480 87.570 ;
        RECT 108.200 86.845 109.200 87.015 ;
        RECT 110.080 86.845 111.080 87.015 ;
        RECT 111.960 86.845 112.960 87.015 ;
        RECT 113.840 86.845 114.840 87.015 ;
        RECT 115.720 86.845 116.720 87.015 ;
        RECT 117.600 86.845 118.600 87.015 ;
        RECT 104.230 86.600 104.730 86.770 ;
        RECT 105.630 86.600 106.130 86.770 ;
        RECT 104.230 86.035 104.730 86.205 ;
        RECT 105.630 86.035 106.130 86.205 ;
        RECT 100.890 84.790 102.540 84.960 ;
        RECT 85.540 82.205 86.540 82.375 ;
        RECT 87.420 82.205 88.420 82.375 ;
        RECT 89.300 82.205 90.300 82.375 ;
        RECT 91.180 82.205 92.180 82.375 ;
        RECT 93.060 82.205 94.060 82.375 ;
        RECT 94.940 82.205 95.940 82.375 ;
        RECT 85.540 81.665 86.540 81.835 ;
        RECT 87.420 81.665 88.420 81.835 ;
        RECT 89.300 81.665 90.300 81.835 ;
        RECT 91.180 81.665 92.180 81.835 ;
        RECT 93.060 81.665 94.060 81.835 ;
        RECT 94.940 81.665 95.940 81.835 ;
        RECT 85.310 77.410 85.480 81.450 ;
        RECT 86.600 77.410 86.770 81.450 ;
        RECT 87.190 77.410 87.360 81.450 ;
        RECT 88.480 77.410 88.650 81.450 ;
        RECT 89.070 77.410 89.240 81.450 ;
        RECT 92.240 77.410 92.410 81.450 ;
        RECT 94.120 77.410 94.290 81.450 ;
        RECT 96.000 77.410 96.170 81.450 ;
        RECT 78.230 77.000 79.880 77.170 ;
        RECT 85.540 77.025 86.540 77.195 ;
        RECT 87.420 77.025 88.420 77.195 ;
        RECT 89.300 77.025 90.300 77.195 ;
        RECT 91.180 77.025 92.180 77.195 ;
        RECT 93.060 77.025 94.060 77.195 ;
        RECT 94.940 77.025 95.940 77.195 ;
        RECT 96.710 76.430 97.060 78.590 ;
        RECT 97.540 76.430 97.890 78.590 ;
        RECT 98.370 76.430 98.720 78.590 ;
        RECT 99.200 76.430 99.550 78.590 ;
        RECT 100.890 77.170 101.060 84.790 ;
        RECT 101.540 82.150 101.890 84.310 ;
        RECT 101.540 77.650 101.890 79.810 ;
        RECT 102.370 77.170 102.540 84.790 ;
        RECT 104.000 84.780 104.170 85.820 ;
        RECT 105.400 84.780 105.570 85.820 ;
        RECT 104.230 84.395 104.730 84.565 ;
        RECT 105.630 84.395 106.130 84.565 ;
        RECT 107.970 82.590 108.140 86.630 ;
        RECT 109.260 82.590 109.430 86.630 ;
        RECT 109.850 82.590 110.020 86.630 ;
        RECT 111.140 82.590 111.310 86.630 ;
        RECT 111.730 82.590 111.900 86.630 ;
        RECT 114.900 82.590 115.070 86.630 ;
        RECT 116.780 82.590 116.950 86.630 ;
        RECT 118.660 82.590 118.830 86.630 ;
        RECT 119.370 84.680 119.720 86.840 ;
        RECT 120.200 84.680 120.550 86.840 ;
        RECT 121.030 84.680 121.380 86.840 ;
        RECT 123.550 84.960 123.720 92.580 ;
        RECT 124.200 89.940 124.550 92.100 ;
        RECT 124.200 85.440 124.550 87.600 ;
        RECT 125.030 84.960 125.200 92.580 ;
        RECT 123.550 84.790 125.200 84.960 ;
        RECT 108.200 82.205 109.200 82.375 ;
        RECT 110.080 82.205 111.080 82.375 ;
        RECT 111.960 82.205 112.960 82.375 ;
        RECT 113.840 82.205 114.840 82.375 ;
        RECT 115.720 82.205 116.720 82.375 ;
        RECT 117.600 82.205 118.600 82.375 ;
        RECT 108.200 81.665 109.200 81.835 ;
        RECT 110.080 81.665 111.080 81.835 ;
        RECT 111.960 81.665 112.960 81.835 ;
        RECT 113.840 81.665 114.840 81.835 ;
        RECT 115.720 81.665 116.720 81.835 ;
        RECT 117.600 81.665 118.600 81.835 ;
        RECT 107.970 77.410 108.140 81.450 ;
        RECT 109.260 77.410 109.430 81.450 ;
        RECT 109.850 77.410 110.020 81.450 ;
        RECT 111.140 77.410 111.310 81.450 ;
        RECT 111.730 77.410 111.900 81.450 ;
        RECT 114.900 77.410 115.070 81.450 ;
        RECT 116.780 77.410 116.950 81.450 ;
        RECT 118.660 77.410 118.830 81.450 ;
        RECT 100.890 77.000 102.540 77.170 ;
        RECT 108.200 77.025 109.200 77.195 ;
        RECT 110.080 77.025 111.080 77.195 ;
        RECT 111.960 77.025 112.960 77.195 ;
        RECT 113.840 77.025 114.840 77.195 ;
        RECT 115.720 77.025 116.720 77.195 ;
        RECT 117.600 77.025 118.600 77.195 ;
        RECT 119.370 76.430 119.720 78.590 ;
        RECT 120.200 76.430 120.550 78.590 ;
        RECT 121.030 76.430 121.380 78.590 ;
        RECT 121.860 76.430 122.210 78.590 ;
        RECT 123.550 77.170 123.720 84.790 ;
        RECT 124.200 82.150 124.550 84.310 ;
        RECT 124.200 77.650 124.550 79.810 ;
        RECT 125.030 77.170 125.200 84.790 ;
        RECT 123.550 77.000 125.200 77.170 ;
        RECT 40.220 75.700 41.220 75.870 ;
        RECT 42.100 75.700 43.100 75.870 ;
        RECT 43.980 75.700 44.980 75.870 ;
        RECT 45.860 75.700 46.860 75.870 ;
        RECT 47.740 75.700 48.740 75.870 ;
        RECT 49.620 75.700 50.620 75.870 ;
        RECT 51.500 75.700 52.500 75.870 ;
        RECT 62.880 75.700 63.880 75.870 ;
        RECT 64.760 75.700 65.760 75.870 ;
        RECT 66.640 75.700 67.640 75.870 ;
        RECT 68.520 75.700 69.520 75.870 ;
        RECT 70.400 75.700 71.400 75.870 ;
        RECT 72.280 75.700 73.280 75.870 ;
        RECT 74.160 75.700 75.160 75.870 ;
        RECT 85.540 75.700 86.540 75.870 ;
        RECT 87.420 75.700 88.420 75.870 ;
        RECT 89.300 75.700 90.300 75.870 ;
        RECT 91.180 75.700 92.180 75.870 ;
        RECT 93.060 75.700 94.060 75.870 ;
        RECT 94.940 75.700 95.940 75.870 ;
        RECT 96.820 75.700 97.820 75.870 ;
        RECT 108.200 75.700 109.200 75.870 ;
        RECT 110.080 75.700 111.080 75.870 ;
        RECT 111.960 75.700 112.960 75.870 ;
        RECT 113.840 75.700 114.840 75.870 ;
        RECT 115.720 75.700 116.720 75.870 ;
        RECT 117.600 75.700 118.600 75.870 ;
        RECT 119.480 75.700 120.480 75.870 ;
        RECT 39.990 73.490 40.160 75.530 ;
        RECT 43.160 73.490 43.330 75.530 ;
        RECT 43.750 73.490 43.920 75.530 ;
        RECT 45.040 73.490 45.210 75.530 ;
        RECT 45.630 73.490 45.800 75.530 ;
        RECT 46.920 73.490 47.090 75.530 ;
        RECT 48.800 73.490 48.970 75.530 ;
        RECT 50.680 73.490 50.850 75.530 ;
        RECT 52.560 73.490 52.730 75.530 ;
        RECT 55.570 75.240 57.220 75.410 ;
        RECT 40.220 73.150 41.220 73.320 ;
        RECT 42.100 73.150 43.100 73.320 ;
        RECT 43.980 73.150 44.980 73.320 ;
        RECT 45.860 73.150 46.860 73.320 ;
        RECT 47.740 73.150 48.740 73.320 ;
        RECT 49.620 73.150 50.620 73.320 ;
        RECT 51.500 73.150 52.500 73.320 ;
        RECT 40.220 72.610 41.220 72.780 ;
        RECT 42.100 72.610 43.100 72.780 ;
        RECT 43.980 72.610 44.980 72.780 ;
        RECT 45.860 72.610 46.860 72.780 ;
        RECT 47.740 72.610 48.740 72.780 ;
        RECT 49.620 72.610 50.620 72.780 ;
        RECT 51.500 72.610 52.500 72.780 ;
        RECT 36.250 70.310 36.750 70.480 ;
        RECT 37.650 70.310 38.150 70.480 ;
        RECT 39.990 70.400 40.160 72.440 ;
        RECT 43.160 70.400 43.330 72.440 ;
        RECT 43.750 70.400 43.920 72.440 ;
        RECT 45.040 70.400 45.210 72.440 ;
        RECT 45.630 70.400 45.800 72.440 ;
        RECT 46.920 70.400 47.090 72.440 ;
        RECT 48.800 70.400 48.970 72.440 ;
        RECT 50.680 70.400 50.850 72.440 ;
        RECT 52.560 70.400 52.730 72.440 ;
        RECT 36.020 69.600 36.190 70.140 ;
        RECT 37.420 69.600 37.590 70.140 ;
        RECT 40.220 70.060 41.220 70.230 ;
        RECT 42.100 70.060 43.100 70.230 ;
        RECT 43.980 70.060 44.980 70.230 ;
        RECT 45.860 70.060 46.860 70.230 ;
        RECT 47.740 70.060 48.740 70.230 ;
        RECT 49.620 70.060 50.620 70.230 ;
        RECT 51.500 70.060 52.500 70.230 ;
        RECT 40.220 69.505 41.220 69.675 ;
        RECT 42.100 69.505 43.100 69.675 ;
        RECT 43.980 69.505 44.980 69.675 ;
        RECT 45.860 69.505 46.860 69.675 ;
        RECT 47.740 69.505 48.740 69.675 ;
        RECT 49.620 69.505 50.620 69.675 ;
        RECT 36.250 69.260 36.750 69.430 ;
        RECT 37.650 69.260 38.150 69.430 ;
        RECT 36.250 68.695 36.750 68.865 ;
        RECT 37.650 68.695 38.150 68.865 ;
        RECT 36.020 67.440 36.190 68.480 ;
        RECT 37.420 67.440 37.590 68.480 ;
        RECT 36.250 67.055 36.750 67.225 ;
        RECT 37.650 67.055 38.150 67.225 ;
        RECT 39.990 65.250 40.160 69.290 ;
        RECT 41.280 65.250 41.450 69.290 ;
        RECT 41.870 65.250 42.040 69.290 ;
        RECT 43.160 65.250 43.330 69.290 ;
        RECT 43.750 65.250 43.920 69.290 ;
        RECT 46.920 65.250 47.090 69.290 ;
        RECT 48.800 65.250 48.970 69.290 ;
        RECT 50.680 65.250 50.850 69.290 ;
        RECT 51.390 67.340 51.740 69.500 ;
        RECT 52.220 67.340 52.570 69.500 ;
        RECT 53.050 67.340 53.400 69.500 ;
        RECT 55.570 67.620 55.740 75.240 ;
        RECT 56.220 72.600 56.570 74.760 ;
        RECT 56.220 68.100 56.570 70.260 ;
        RECT 57.050 67.620 57.220 75.240 ;
        RECT 62.650 73.490 62.820 75.530 ;
        RECT 65.820 73.490 65.990 75.530 ;
        RECT 66.410 73.490 66.580 75.530 ;
        RECT 67.700 73.490 67.870 75.530 ;
        RECT 68.290 73.490 68.460 75.530 ;
        RECT 69.580 73.490 69.750 75.530 ;
        RECT 71.460 73.490 71.630 75.530 ;
        RECT 73.340 73.490 73.510 75.530 ;
        RECT 75.220 73.490 75.390 75.530 ;
        RECT 78.230 75.240 79.880 75.410 ;
        RECT 62.880 73.150 63.880 73.320 ;
        RECT 64.760 73.150 65.760 73.320 ;
        RECT 66.640 73.150 67.640 73.320 ;
        RECT 68.520 73.150 69.520 73.320 ;
        RECT 70.400 73.150 71.400 73.320 ;
        RECT 72.280 73.150 73.280 73.320 ;
        RECT 74.160 73.150 75.160 73.320 ;
        RECT 62.880 72.610 63.880 72.780 ;
        RECT 64.760 72.610 65.760 72.780 ;
        RECT 66.640 72.610 67.640 72.780 ;
        RECT 68.520 72.610 69.520 72.780 ;
        RECT 70.400 72.610 71.400 72.780 ;
        RECT 72.280 72.610 73.280 72.780 ;
        RECT 74.160 72.610 75.160 72.780 ;
        RECT 58.910 70.310 59.410 70.480 ;
        RECT 60.310 70.310 60.810 70.480 ;
        RECT 62.650 70.400 62.820 72.440 ;
        RECT 65.820 70.400 65.990 72.440 ;
        RECT 66.410 70.400 66.580 72.440 ;
        RECT 67.700 70.400 67.870 72.440 ;
        RECT 68.290 70.400 68.460 72.440 ;
        RECT 69.580 70.400 69.750 72.440 ;
        RECT 71.460 70.400 71.630 72.440 ;
        RECT 73.340 70.400 73.510 72.440 ;
        RECT 75.220 70.400 75.390 72.440 ;
        RECT 58.680 69.600 58.850 70.140 ;
        RECT 60.080 69.600 60.250 70.140 ;
        RECT 62.880 70.060 63.880 70.230 ;
        RECT 64.760 70.060 65.760 70.230 ;
        RECT 66.640 70.060 67.640 70.230 ;
        RECT 68.520 70.060 69.520 70.230 ;
        RECT 70.400 70.060 71.400 70.230 ;
        RECT 72.280 70.060 73.280 70.230 ;
        RECT 74.160 70.060 75.160 70.230 ;
        RECT 62.880 69.505 63.880 69.675 ;
        RECT 64.760 69.505 65.760 69.675 ;
        RECT 66.640 69.505 67.640 69.675 ;
        RECT 68.520 69.505 69.520 69.675 ;
        RECT 70.400 69.505 71.400 69.675 ;
        RECT 72.280 69.505 73.280 69.675 ;
        RECT 58.910 69.260 59.410 69.430 ;
        RECT 60.310 69.260 60.810 69.430 ;
        RECT 58.910 68.695 59.410 68.865 ;
        RECT 60.310 68.695 60.810 68.865 ;
        RECT 55.570 67.450 57.220 67.620 ;
        RECT 40.220 64.865 41.220 65.035 ;
        RECT 42.100 64.865 43.100 65.035 ;
        RECT 43.980 64.865 44.980 65.035 ;
        RECT 45.860 64.865 46.860 65.035 ;
        RECT 47.740 64.865 48.740 65.035 ;
        RECT 49.620 64.865 50.620 65.035 ;
        RECT 40.220 64.325 41.220 64.495 ;
        RECT 42.100 64.325 43.100 64.495 ;
        RECT 43.980 64.325 44.980 64.495 ;
        RECT 45.860 64.325 46.860 64.495 ;
        RECT 47.740 64.325 48.740 64.495 ;
        RECT 49.620 64.325 50.620 64.495 ;
        RECT 39.990 60.070 40.160 64.110 ;
        RECT 41.280 60.070 41.450 64.110 ;
        RECT 41.870 60.070 42.040 64.110 ;
        RECT 43.160 60.070 43.330 64.110 ;
        RECT 43.750 60.070 43.920 64.110 ;
        RECT 46.920 60.070 47.090 64.110 ;
        RECT 48.800 60.070 48.970 64.110 ;
        RECT 50.680 60.070 50.850 64.110 ;
        RECT 40.220 59.685 41.220 59.855 ;
        RECT 42.100 59.685 43.100 59.855 ;
        RECT 43.980 59.685 44.980 59.855 ;
        RECT 45.860 59.685 46.860 59.855 ;
        RECT 47.740 59.685 48.740 59.855 ;
        RECT 49.620 59.685 50.620 59.855 ;
        RECT 51.390 59.090 51.740 61.250 ;
        RECT 52.220 59.090 52.570 61.250 ;
        RECT 53.050 59.090 53.400 61.250 ;
        RECT 53.880 59.090 54.230 61.250 ;
        RECT 55.570 59.830 55.740 67.450 ;
        RECT 56.220 64.810 56.570 66.970 ;
        RECT 56.220 60.310 56.570 62.470 ;
        RECT 57.050 59.830 57.220 67.450 ;
        RECT 58.680 67.440 58.850 68.480 ;
        RECT 60.080 67.440 60.250 68.480 ;
        RECT 58.910 67.055 59.410 67.225 ;
        RECT 60.310 67.055 60.810 67.225 ;
        RECT 62.650 65.250 62.820 69.290 ;
        RECT 63.940 65.250 64.110 69.290 ;
        RECT 64.530 65.250 64.700 69.290 ;
        RECT 65.820 65.250 65.990 69.290 ;
        RECT 66.410 65.250 66.580 69.290 ;
        RECT 69.580 65.250 69.750 69.290 ;
        RECT 71.460 65.250 71.630 69.290 ;
        RECT 73.340 65.250 73.510 69.290 ;
        RECT 74.050 67.340 74.400 69.500 ;
        RECT 74.880 67.340 75.230 69.500 ;
        RECT 75.710 67.340 76.060 69.500 ;
        RECT 78.230 67.620 78.400 75.240 ;
        RECT 78.880 72.600 79.230 74.760 ;
        RECT 78.880 68.100 79.230 70.260 ;
        RECT 79.710 67.620 79.880 75.240 ;
        RECT 85.310 73.490 85.480 75.530 ;
        RECT 88.480 73.490 88.650 75.530 ;
        RECT 89.070 73.490 89.240 75.530 ;
        RECT 90.360 73.490 90.530 75.530 ;
        RECT 90.950 73.490 91.120 75.530 ;
        RECT 92.240 73.490 92.410 75.530 ;
        RECT 94.120 73.490 94.290 75.530 ;
        RECT 96.000 73.490 96.170 75.530 ;
        RECT 97.880 73.490 98.050 75.530 ;
        RECT 100.890 75.240 102.540 75.410 ;
        RECT 85.540 73.150 86.540 73.320 ;
        RECT 87.420 73.150 88.420 73.320 ;
        RECT 89.300 73.150 90.300 73.320 ;
        RECT 91.180 73.150 92.180 73.320 ;
        RECT 93.060 73.150 94.060 73.320 ;
        RECT 94.940 73.150 95.940 73.320 ;
        RECT 96.820 73.150 97.820 73.320 ;
        RECT 85.540 72.610 86.540 72.780 ;
        RECT 87.420 72.610 88.420 72.780 ;
        RECT 89.300 72.610 90.300 72.780 ;
        RECT 91.180 72.610 92.180 72.780 ;
        RECT 93.060 72.610 94.060 72.780 ;
        RECT 94.940 72.610 95.940 72.780 ;
        RECT 96.820 72.610 97.820 72.780 ;
        RECT 81.570 70.310 82.070 70.480 ;
        RECT 82.970 70.310 83.470 70.480 ;
        RECT 85.310 70.400 85.480 72.440 ;
        RECT 88.480 70.400 88.650 72.440 ;
        RECT 89.070 70.400 89.240 72.440 ;
        RECT 90.360 70.400 90.530 72.440 ;
        RECT 90.950 70.400 91.120 72.440 ;
        RECT 92.240 70.400 92.410 72.440 ;
        RECT 94.120 70.400 94.290 72.440 ;
        RECT 96.000 70.400 96.170 72.440 ;
        RECT 97.880 70.400 98.050 72.440 ;
        RECT 81.340 69.600 81.510 70.140 ;
        RECT 82.740 69.600 82.910 70.140 ;
        RECT 85.540 70.060 86.540 70.230 ;
        RECT 87.420 70.060 88.420 70.230 ;
        RECT 89.300 70.060 90.300 70.230 ;
        RECT 91.180 70.060 92.180 70.230 ;
        RECT 93.060 70.060 94.060 70.230 ;
        RECT 94.940 70.060 95.940 70.230 ;
        RECT 96.820 70.060 97.820 70.230 ;
        RECT 85.540 69.505 86.540 69.675 ;
        RECT 87.420 69.505 88.420 69.675 ;
        RECT 89.300 69.505 90.300 69.675 ;
        RECT 91.180 69.505 92.180 69.675 ;
        RECT 93.060 69.505 94.060 69.675 ;
        RECT 94.940 69.505 95.940 69.675 ;
        RECT 81.570 69.260 82.070 69.430 ;
        RECT 82.970 69.260 83.470 69.430 ;
        RECT 81.570 68.695 82.070 68.865 ;
        RECT 82.970 68.695 83.470 68.865 ;
        RECT 78.230 67.450 79.880 67.620 ;
        RECT 62.880 64.865 63.880 65.035 ;
        RECT 64.760 64.865 65.760 65.035 ;
        RECT 66.640 64.865 67.640 65.035 ;
        RECT 68.520 64.865 69.520 65.035 ;
        RECT 70.400 64.865 71.400 65.035 ;
        RECT 72.280 64.865 73.280 65.035 ;
        RECT 62.880 64.325 63.880 64.495 ;
        RECT 64.760 64.325 65.760 64.495 ;
        RECT 66.640 64.325 67.640 64.495 ;
        RECT 68.520 64.325 69.520 64.495 ;
        RECT 70.400 64.325 71.400 64.495 ;
        RECT 72.280 64.325 73.280 64.495 ;
        RECT 62.650 60.070 62.820 64.110 ;
        RECT 63.940 60.070 64.110 64.110 ;
        RECT 64.530 60.070 64.700 64.110 ;
        RECT 65.820 60.070 65.990 64.110 ;
        RECT 66.410 60.070 66.580 64.110 ;
        RECT 69.580 60.070 69.750 64.110 ;
        RECT 71.460 60.070 71.630 64.110 ;
        RECT 73.340 60.070 73.510 64.110 ;
        RECT 55.570 59.660 57.220 59.830 ;
        RECT 62.880 59.685 63.880 59.855 ;
        RECT 64.760 59.685 65.760 59.855 ;
        RECT 66.640 59.685 67.640 59.855 ;
        RECT 68.520 59.685 69.520 59.855 ;
        RECT 70.400 59.685 71.400 59.855 ;
        RECT 72.280 59.685 73.280 59.855 ;
        RECT 74.050 59.090 74.400 61.250 ;
        RECT 74.880 59.090 75.230 61.250 ;
        RECT 75.710 59.090 76.060 61.250 ;
        RECT 76.540 59.090 76.890 61.250 ;
        RECT 78.230 59.830 78.400 67.450 ;
        RECT 78.880 64.810 79.230 66.970 ;
        RECT 78.880 60.310 79.230 62.470 ;
        RECT 79.710 59.830 79.880 67.450 ;
        RECT 81.340 67.440 81.510 68.480 ;
        RECT 82.740 67.440 82.910 68.480 ;
        RECT 81.570 67.055 82.070 67.225 ;
        RECT 82.970 67.055 83.470 67.225 ;
        RECT 85.310 65.250 85.480 69.290 ;
        RECT 86.600 65.250 86.770 69.290 ;
        RECT 87.190 65.250 87.360 69.290 ;
        RECT 88.480 65.250 88.650 69.290 ;
        RECT 89.070 65.250 89.240 69.290 ;
        RECT 92.240 65.250 92.410 69.290 ;
        RECT 94.120 65.250 94.290 69.290 ;
        RECT 96.000 65.250 96.170 69.290 ;
        RECT 96.710 67.340 97.060 69.500 ;
        RECT 97.540 67.340 97.890 69.500 ;
        RECT 98.370 67.340 98.720 69.500 ;
        RECT 100.890 67.620 101.060 75.240 ;
        RECT 101.540 72.600 101.890 74.760 ;
        RECT 101.540 68.100 101.890 70.260 ;
        RECT 102.370 67.620 102.540 75.240 ;
        RECT 107.970 73.490 108.140 75.530 ;
        RECT 111.140 73.490 111.310 75.530 ;
        RECT 111.730 73.490 111.900 75.530 ;
        RECT 113.020 73.490 113.190 75.530 ;
        RECT 113.610 73.490 113.780 75.530 ;
        RECT 114.900 73.490 115.070 75.530 ;
        RECT 116.780 73.490 116.950 75.530 ;
        RECT 118.660 73.490 118.830 75.530 ;
        RECT 120.540 73.490 120.710 75.530 ;
        RECT 123.550 75.240 125.200 75.410 ;
        RECT 108.200 73.150 109.200 73.320 ;
        RECT 110.080 73.150 111.080 73.320 ;
        RECT 111.960 73.150 112.960 73.320 ;
        RECT 113.840 73.150 114.840 73.320 ;
        RECT 115.720 73.150 116.720 73.320 ;
        RECT 117.600 73.150 118.600 73.320 ;
        RECT 119.480 73.150 120.480 73.320 ;
        RECT 108.200 72.610 109.200 72.780 ;
        RECT 110.080 72.610 111.080 72.780 ;
        RECT 111.960 72.610 112.960 72.780 ;
        RECT 113.840 72.610 114.840 72.780 ;
        RECT 115.720 72.610 116.720 72.780 ;
        RECT 117.600 72.610 118.600 72.780 ;
        RECT 119.480 72.610 120.480 72.780 ;
        RECT 104.230 70.310 104.730 70.480 ;
        RECT 105.630 70.310 106.130 70.480 ;
        RECT 107.970 70.400 108.140 72.440 ;
        RECT 111.140 70.400 111.310 72.440 ;
        RECT 111.730 70.400 111.900 72.440 ;
        RECT 113.020 70.400 113.190 72.440 ;
        RECT 113.610 70.400 113.780 72.440 ;
        RECT 114.900 70.400 115.070 72.440 ;
        RECT 116.780 70.400 116.950 72.440 ;
        RECT 118.660 70.400 118.830 72.440 ;
        RECT 120.540 70.400 120.710 72.440 ;
        RECT 104.000 69.600 104.170 70.140 ;
        RECT 105.400 69.600 105.570 70.140 ;
        RECT 108.200 70.060 109.200 70.230 ;
        RECT 110.080 70.060 111.080 70.230 ;
        RECT 111.960 70.060 112.960 70.230 ;
        RECT 113.840 70.060 114.840 70.230 ;
        RECT 115.720 70.060 116.720 70.230 ;
        RECT 117.600 70.060 118.600 70.230 ;
        RECT 119.480 70.060 120.480 70.230 ;
        RECT 108.200 69.505 109.200 69.675 ;
        RECT 110.080 69.505 111.080 69.675 ;
        RECT 111.960 69.505 112.960 69.675 ;
        RECT 113.840 69.505 114.840 69.675 ;
        RECT 115.720 69.505 116.720 69.675 ;
        RECT 117.600 69.505 118.600 69.675 ;
        RECT 104.230 69.260 104.730 69.430 ;
        RECT 105.630 69.260 106.130 69.430 ;
        RECT 104.230 68.695 104.730 68.865 ;
        RECT 105.630 68.695 106.130 68.865 ;
        RECT 100.890 67.450 102.540 67.620 ;
        RECT 85.540 64.865 86.540 65.035 ;
        RECT 87.420 64.865 88.420 65.035 ;
        RECT 89.300 64.865 90.300 65.035 ;
        RECT 91.180 64.865 92.180 65.035 ;
        RECT 93.060 64.865 94.060 65.035 ;
        RECT 94.940 64.865 95.940 65.035 ;
        RECT 85.540 64.325 86.540 64.495 ;
        RECT 87.420 64.325 88.420 64.495 ;
        RECT 89.300 64.325 90.300 64.495 ;
        RECT 91.180 64.325 92.180 64.495 ;
        RECT 93.060 64.325 94.060 64.495 ;
        RECT 94.940 64.325 95.940 64.495 ;
        RECT 85.310 60.070 85.480 64.110 ;
        RECT 86.600 60.070 86.770 64.110 ;
        RECT 87.190 60.070 87.360 64.110 ;
        RECT 88.480 60.070 88.650 64.110 ;
        RECT 89.070 60.070 89.240 64.110 ;
        RECT 92.240 60.070 92.410 64.110 ;
        RECT 94.120 60.070 94.290 64.110 ;
        RECT 96.000 60.070 96.170 64.110 ;
        RECT 78.230 59.660 79.880 59.830 ;
        RECT 85.540 59.685 86.540 59.855 ;
        RECT 87.420 59.685 88.420 59.855 ;
        RECT 89.300 59.685 90.300 59.855 ;
        RECT 91.180 59.685 92.180 59.855 ;
        RECT 93.060 59.685 94.060 59.855 ;
        RECT 94.940 59.685 95.940 59.855 ;
        RECT 96.710 59.090 97.060 61.250 ;
        RECT 97.540 59.090 97.890 61.250 ;
        RECT 98.370 59.090 98.720 61.250 ;
        RECT 99.200 59.090 99.550 61.250 ;
        RECT 100.890 59.830 101.060 67.450 ;
        RECT 101.540 64.810 101.890 66.970 ;
        RECT 101.540 60.310 101.890 62.470 ;
        RECT 102.370 59.830 102.540 67.450 ;
        RECT 104.000 67.440 104.170 68.480 ;
        RECT 105.400 67.440 105.570 68.480 ;
        RECT 104.230 67.055 104.730 67.225 ;
        RECT 105.630 67.055 106.130 67.225 ;
        RECT 107.970 65.250 108.140 69.290 ;
        RECT 109.260 65.250 109.430 69.290 ;
        RECT 109.850 65.250 110.020 69.290 ;
        RECT 111.140 65.250 111.310 69.290 ;
        RECT 111.730 65.250 111.900 69.290 ;
        RECT 114.900 65.250 115.070 69.290 ;
        RECT 116.780 65.250 116.950 69.290 ;
        RECT 118.660 65.250 118.830 69.290 ;
        RECT 119.370 67.340 119.720 69.500 ;
        RECT 120.200 67.340 120.550 69.500 ;
        RECT 121.030 67.340 121.380 69.500 ;
        RECT 123.550 67.620 123.720 75.240 ;
        RECT 124.200 72.600 124.550 74.760 ;
        RECT 124.200 68.100 124.550 70.260 ;
        RECT 125.030 67.620 125.200 75.240 ;
        RECT 123.550 67.450 125.200 67.620 ;
        RECT 108.200 64.865 109.200 65.035 ;
        RECT 110.080 64.865 111.080 65.035 ;
        RECT 111.960 64.865 112.960 65.035 ;
        RECT 113.840 64.865 114.840 65.035 ;
        RECT 115.720 64.865 116.720 65.035 ;
        RECT 117.600 64.865 118.600 65.035 ;
        RECT 108.200 64.325 109.200 64.495 ;
        RECT 110.080 64.325 111.080 64.495 ;
        RECT 111.960 64.325 112.960 64.495 ;
        RECT 113.840 64.325 114.840 64.495 ;
        RECT 115.720 64.325 116.720 64.495 ;
        RECT 117.600 64.325 118.600 64.495 ;
        RECT 107.970 60.070 108.140 64.110 ;
        RECT 109.260 60.070 109.430 64.110 ;
        RECT 109.850 60.070 110.020 64.110 ;
        RECT 111.140 60.070 111.310 64.110 ;
        RECT 111.730 60.070 111.900 64.110 ;
        RECT 114.900 60.070 115.070 64.110 ;
        RECT 116.780 60.070 116.950 64.110 ;
        RECT 118.660 60.070 118.830 64.110 ;
        RECT 100.890 59.660 102.540 59.830 ;
        RECT 108.200 59.685 109.200 59.855 ;
        RECT 110.080 59.685 111.080 59.855 ;
        RECT 111.960 59.685 112.960 59.855 ;
        RECT 113.840 59.685 114.840 59.855 ;
        RECT 115.720 59.685 116.720 59.855 ;
        RECT 117.600 59.685 118.600 59.855 ;
        RECT 119.370 59.090 119.720 61.250 ;
        RECT 120.200 59.090 120.550 61.250 ;
        RECT 121.030 59.090 121.380 61.250 ;
        RECT 121.860 59.090 122.210 61.250 ;
        RECT 123.550 59.830 123.720 67.450 ;
        RECT 124.200 64.810 124.550 66.970 ;
        RECT 124.200 60.310 124.550 62.470 ;
        RECT 125.030 59.830 125.200 67.450 ;
        RECT 123.550 59.660 125.200 59.830 ;
        RECT 40.220 57.700 41.220 57.870 ;
        RECT 42.100 57.700 43.100 57.870 ;
        RECT 43.980 57.700 44.980 57.870 ;
        RECT 47.740 57.700 48.740 57.870 ;
        RECT 49.620 57.700 50.620 57.870 ;
        RECT 51.500 57.700 52.500 57.870 ;
        RECT 62.880 57.700 63.880 57.870 ;
        RECT 64.760 57.700 65.760 57.870 ;
        RECT 66.640 57.700 67.640 57.870 ;
        RECT 70.400 57.700 71.400 57.870 ;
        RECT 72.280 57.700 73.280 57.870 ;
        RECT 74.160 57.700 75.160 57.870 ;
        RECT 85.540 57.700 86.540 57.870 ;
        RECT 87.420 57.700 88.420 57.870 ;
        RECT 89.300 57.700 90.300 57.870 ;
        RECT 93.060 57.700 94.060 57.870 ;
        RECT 94.940 57.700 95.940 57.870 ;
        RECT 96.820 57.700 97.820 57.870 ;
        RECT 108.200 57.700 109.200 57.870 ;
        RECT 110.080 57.700 111.080 57.870 ;
        RECT 111.960 57.700 112.960 57.870 ;
        RECT 115.720 57.700 116.720 57.870 ;
        RECT 117.600 57.700 118.600 57.870 ;
        RECT 119.480 57.700 120.480 57.870 ;
        RECT 39.990 55.490 40.160 57.530 ;
        RECT 43.160 55.490 43.330 57.530 ;
        RECT 43.750 55.490 43.920 57.530 ;
        RECT 45.040 55.490 45.210 57.530 ;
        RECT 45.630 55.490 45.800 57.530 ;
        RECT 46.920 55.490 47.090 57.530 ;
        RECT 48.800 55.490 48.970 57.530 ;
        RECT 50.680 55.490 50.850 57.530 ;
        RECT 52.560 55.490 52.730 57.530 ;
        RECT 62.650 55.490 62.820 57.530 ;
        RECT 65.820 55.490 65.990 57.530 ;
        RECT 66.410 55.490 66.580 57.530 ;
        RECT 67.700 55.490 67.870 57.530 ;
        RECT 68.290 55.490 68.460 57.530 ;
        RECT 69.580 55.490 69.750 57.530 ;
        RECT 71.460 55.490 71.630 57.530 ;
        RECT 73.340 55.490 73.510 57.530 ;
        RECT 75.220 55.490 75.390 57.530 ;
        RECT 85.310 55.490 85.480 57.530 ;
        RECT 88.480 55.490 88.650 57.530 ;
        RECT 89.070 55.490 89.240 57.530 ;
        RECT 90.360 55.490 90.530 57.530 ;
        RECT 90.950 55.490 91.120 57.530 ;
        RECT 92.240 55.490 92.410 57.530 ;
        RECT 94.120 55.490 94.290 57.530 ;
        RECT 96.000 55.490 96.170 57.530 ;
        RECT 97.880 55.490 98.050 57.530 ;
        RECT 107.970 55.490 108.140 57.530 ;
        RECT 111.140 55.490 111.310 57.530 ;
        RECT 111.730 55.490 111.900 57.530 ;
        RECT 113.020 55.490 113.190 57.530 ;
        RECT 113.610 55.490 113.780 57.530 ;
        RECT 114.900 55.490 115.070 57.530 ;
        RECT 116.780 55.490 116.950 57.530 ;
        RECT 118.660 55.490 118.830 57.530 ;
        RECT 120.540 55.490 120.710 57.530 ;
        RECT 40.220 55.150 41.220 55.320 ;
        RECT 42.100 55.150 43.100 55.320 ;
        RECT 43.980 55.150 44.980 55.320 ;
        RECT 47.740 55.150 48.740 55.320 ;
        RECT 49.620 55.150 50.620 55.320 ;
        RECT 51.500 55.150 52.500 55.320 ;
        RECT 62.880 55.150 63.880 55.320 ;
        RECT 64.760 55.150 65.760 55.320 ;
        RECT 66.640 55.150 67.640 55.320 ;
        RECT 70.400 55.150 71.400 55.320 ;
        RECT 72.280 55.150 73.280 55.320 ;
        RECT 74.160 55.150 75.160 55.320 ;
        RECT 85.540 55.150 86.540 55.320 ;
        RECT 87.420 55.150 88.420 55.320 ;
        RECT 89.300 55.150 90.300 55.320 ;
        RECT 93.060 55.150 94.060 55.320 ;
        RECT 94.940 55.150 95.940 55.320 ;
        RECT 96.820 55.150 97.820 55.320 ;
        RECT 108.200 55.150 109.200 55.320 ;
        RECT 110.080 55.150 111.080 55.320 ;
        RECT 111.960 55.150 112.960 55.320 ;
        RECT 115.720 55.150 116.720 55.320 ;
        RECT 117.600 55.150 118.600 55.320 ;
        RECT 119.480 55.150 120.480 55.320 ;
        RECT 40.220 54.610 41.220 54.780 ;
        RECT 42.100 54.610 43.100 54.780 ;
        RECT 43.980 54.610 44.980 54.780 ;
        RECT 47.740 54.610 48.740 54.780 ;
        RECT 49.620 54.610 50.620 54.780 ;
        RECT 51.500 54.610 52.500 54.780 ;
        RECT 62.880 54.610 63.880 54.780 ;
        RECT 64.760 54.610 65.760 54.780 ;
        RECT 66.640 54.610 67.640 54.780 ;
        RECT 70.400 54.610 71.400 54.780 ;
        RECT 72.280 54.610 73.280 54.780 ;
        RECT 74.160 54.610 75.160 54.780 ;
        RECT 85.540 54.610 86.540 54.780 ;
        RECT 87.420 54.610 88.420 54.780 ;
        RECT 89.300 54.610 90.300 54.780 ;
        RECT 93.060 54.610 94.060 54.780 ;
        RECT 94.940 54.610 95.940 54.780 ;
        RECT 96.820 54.610 97.820 54.780 ;
        RECT 108.200 54.610 109.200 54.780 ;
        RECT 110.080 54.610 111.080 54.780 ;
        RECT 111.960 54.610 112.960 54.780 ;
        RECT 115.720 54.610 116.720 54.780 ;
        RECT 117.600 54.610 118.600 54.780 ;
        RECT 119.480 54.610 120.480 54.780 ;
        RECT 39.990 52.400 40.160 54.440 ;
        RECT 43.160 52.400 43.330 54.440 ;
        RECT 43.750 52.400 43.920 54.440 ;
        RECT 45.040 52.400 45.210 54.440 ;
        RECT 45.630 52.400 45.800 54.440 ;
        RECT 46.920 52.400 47.090 54.440 ;
        RECT 48.800 52.400 48.970 54.440 ;
        RECT 50.680 52.400 50.850 54.440 ;
        RECT 52.560 52.400 52.730 54.440 ;
        RECT 62.650 52.400 62.820 54.440 ;
        RECT 65.820 52.400 65.990 54.440 ;
        RECT 66.410 52.400 66.580 54.440 ;
        RECT 67.700 52.400 67.870 54.440 ;
        RECT 68.290 52.400 68.460 54.440 ;
        RECT 69.580 52.400 69.750 54.440 ;
        RECT 71.460 52.400 71.630 54.440 ;
        RECT 73.340 52.400 73.510 54.440 ;
        RECT 75.220 52.400 75.390 54.440 ;
        RECT 85.310 52.400 85.480 54.440 ;
        RECT 88.480 52.400 88.650 54.440 ;
        RECT 89.070 52.400 89.240 54.440 ;
        RECT 90.360 52.400 90.530 54.440 ;
        RECT 90.950 52.400 91.120 54.440 ;
        RECT 92.240 52.400 92.410 54.440 ;
        RECT 94.120 52.400 94.290 54.440 ;
        RECT 96.000 52.400 96.170 54.440 ;
        RECT 97.880 52.400 98.050 54.440 ;
        RECT 107.970 52.400 108.140 54.440 ;
        RECT 111.140 52.400 111.310 54.440 ;
        RECT 111.730 52.400 111.900 54.440 ;
        RECT 113.020 52.400 113.190 54.440 ;
        RECT 113.610 52.400 113.780 54.440 ;
        RECT 114.900 52.400 115.070 54.440 ;
        RECT 116.780 52.400 116.950 54.440 ;
        RECT 118.660 52.400 118.830 54.440 ;
        RECT 120.540 52.400 120.710 54.440 ;
        RECT 40.220 52.060 41.220 52.230 ;
        RECT 42.100 52.060 43.100 52.230 ;
        RECT 43.980 52.060 44.980 52.230 ;
        RECT 47.740 52.060 48.740 52.230 ;
        RECT 49.620 52.060 50.620 52.230 ;
        RECT 51.500 52.060 52.500 52.230 ;
        RECT 62.880 52.060 63.880 52.230 ;
        RECT 64.760 52.060 65.760 52.230 ;
        RECT 66.640 52.060 67.640 52.230 ;
        RECT 70.400 52.060 71.400 52.230 ;
        RECT 72.280 52.060 73.280 52.230 ;
        RECT 74.160 52.060 75.160 52.230 ;
        RECT 85.540 52.060 86.540 52.230 ;
        RECT 87.420 52.060 88.420 52.230 ;
        RECT 89.300 52.060 90.300 52.230 ;
        RECT 93.060 52.060 94.060 52.230 ;
        RECT 94.940 52.060 95.940 52.230 ;
        RECT 96.820 52.060 97.820 52.230 ;
        RECT 108.200 52.060 109.200 52.230 ;
        RECT 110.080 52.060 111.080 52.230 ;
        RECT 111.960 52.060 112.960 52.230 ;
        RECT 115.720 52.060 116.720 52.230 ;
        RECT 117.600 52.060 118.600 52.230 ;
        RECT 119.480 52.060 120.480 52.230 ;
        RECT 40.220 51.505 41.220 51.675 ;
        RECT 43.980 51.505 44.980 51.675 ;
        RECT 45.860 51.505 46.860 51.675 ;
        RECT 47.740 51.505 48.740 51.675 ;
        RECT 49.620 51.505 50.620 51.675 ;
        RECT 62.880 51.505 63.880 51.675 ;
        RECT 66.640 51.505 67.640 51.675 ;
        RECT 68.520 51.505 69.520 51.675 ;
        RECT 70.400 51.505 71.400 51.675 ;
        RECT 72.280 51.505 73.280 51.675 ;
        RECT 85.540 51.505 86.540 51.675 ;
        RECT 89.300 51.505 90.300 51.675 ;
        RECT 91.180 51.505 92.180 51.675 ;
        RECT 93.060 51.505 94.060 51.675 ;
        RECT 94.940 51.505 95.940 51.675 ;
        RECT 108.200 51.505 109.200 51.675 ;
        RECT 111.960 51.505 112.960 51.675 ;
        RECT 113.840 51.505 114.840 51.675 ;
        RECT 115.720 51.505 116.720 51.675 ;
        RECT 117.600 51.505 118.600 51.675 ;
        RECT 39.990 47.250 40.160 51.290 ;
        RECT 41.280 47.250 41.450 51.290 ;
        RECT 41.870 47.250 42.040 51.290 ;
        RECT 43.160 47.250 43.330 51.290 ;
        RECT 43.750 47.250 43.920 51.290 ;
        RECT 46.920 47.250 47.090 51.290 ;
        RECT 48.800 47.250 48.970 51.290 ;
        RECT 50.680 47.250 50.850 51.290 ;
        RECT 51.390 49.340 51.740 51.500 ;
        RECT 52.220 49.340 52.570 51.500 ;
        RECT 53.050 49.340 53.400 51.500 ;
        RECT 62.650 47.250 62.820 51.290 ;
        RECT 63.940 47.250 64.110 51.290 ;
        RECT 64.530 47.250 64.700 51.290 ;
        RECT 65.820 47.250 65.990 51.290 ;
        RECT 66.410 47.250 66.580 51.290 ;
        RECT 69.580 47.250 69.750 51.290 ;
        RECT 71.460 47.250 71.630 51.290 ;
        RECT 73.340 47.250 73.510 51.290 ;
        RECT 74.050 49.340 74.400 51.500 ;
        RECT 74.880 49.340 75.230 51.500 ;
        RECT 75.710 49.340 76.060 51.500 ;
        RECT 85.310 47.250 85.480 51.290 ;
        RECT 86.600 47.250 86.770 51.290 ;
        RECT 87.190 47.250 87.360 51.290 ;
        RECT 88.480 47.250 88.650 51.290 ;
        RECT 89.070 47.250 89.240 51.290 ;
        RECT 92.240 47.250 92.410 51.290 ;
        RECT 94.120 47.250 94.290 51.290 ;
        RECT 96.000 47.250 96.170 51.290 ;
        RECT 96.710 49.340 97.060 51.500 ;
        RECT 97.540 49.340 97.890 51.500 ;
        RECT 98.370 49.340 98.720 51.500 ;
        RECT 107.970 47.250 108.140 51.290 ;
        RECT 109.260 47.250 109.430 51.290 ;
        RECT 109.850 47.250 110.020 51.290 ;
        RECT 111.140 47.250 111.310 51.290 ;
        RECT 111.730 47.250 111.900 51.290 ;
        RECT 114.900 47.250 115.070 51.290 ;
        RECT 116.780 47.250 116.950 51.290 ;
        RECT 118.660 47.250 118.830 51.290 ;
        RECT 119.370 49.340 119.720 51.500 ;
        RECT 120.200 49.340 120.550 51.500 ;
        RECT 121.030 49.340 121.380 51.500 ;
        RECT 40.220 46.865 41.220 47.035 ;
        RECT 43.980 46.865 44.980 47.035 ;
        RECT 45.860 46.865 46.860 47.035 ;
        RECT 47.740 46.865 48.740 47.035 ;
        RECT 49.620 46.865 50.620 47.035 ;
        RECT 62.880 46.865 63.880 47.035 ;
        RECT 66.640 46.865 67.640 47.035 ;
        RECT 68.520 46.865 69.520 47.035 ;
        RECT 70.400 46.865 71.400 47.035 ;
        RECT 72.280 46.865 73.280 47.035 ;
        RECT 85.540 46.865 86.540 47.035 ;
        RECT 89.300 46.865 90.300 47.035 ;
        RECT 91.180 46.865 92.180 47.035 ;
        RECT 93.060 46.865 94.060 47.035 ;
        RECT 94.940 46.865 95.940 47.035 ;
        RECT 108.200 46.865 109.200 47.035 ;
        RECT 111.960 46.865 112.960 47.035 ;
        RECT 113.840 46.865 114.840 47.035 ;
        RECT 115.720 46.865 116.720 47.035 ;
        RECT 117.600 46.865 118.600 47.035 ;
        RECT 40.220 46.325 41.220 46.495 ;
        RECT 43.980 46.325 44.980 46.495 ;
        RECT 45.860 46.325 46.860 46.495 ;
        RECT 47.740 46.325 48.740 46.495 ;
        RECT 49.620 46.325 50.620 46.495 ;
        RECT 62.880 46.325 63.880 46.495 ;
        RECT 66.640 46.325 67.640 46.495 ;
        RECT 68.520 46.325 69.520 46.495 ;
        RECT 70.400 46.325 71.400 46.495 ;
        RECT 72.280 46.325 73.280 46.495 ;
        RECT 85.540 46.325 86.540 46.495 ;
        RECT 89.300 46.325 90.300 46.495 ;
        RECT 91.180 46.325 92.180 46.495 ;
        RECT 93.060 46.325 94.060 46.495 ;
        RECT 94.940 46.325 95.940 46.495 ;
        RECT 108.200 46.325 109.200 46.495 ;
        RECT 111.960 46.325 112.960 46.495 ;
        RECT 113.840 46.325 114.840 46.495 ;
        RECT 115.720 46.325 116.720 46.495 ;
        RECT 117.600 46.325 118.600 46.495 ;
        RECT 39.990 42.070 40.160 46.110 ;
        RECT 41.280 42.070 41.450 46.110 ;
        RECT 41.870 42.070 42.040 46.110 ;
        RECT 43.160 42.070 43.330 46.110 ;
        RECT 43.750 42.070 43.920 46.110 ;
        RECT 46.920 42.070 47.090 46.110 ;
        RECT 48.800 42.070 48.970 46.110 ;
        RECT 50.680 42.070 50.850 46.110 ;
        RECT 40.220 41.685 41.220 41.855 ;
        RECT 43.980 41.685 44.980 41.855 ;
        RECT 45.860 41.685 46.860 41.855 ;
        RECT 47.740 41.685 48.740 41.855 ;
        RECT 49.620 41.685 50.620 41.855 ;
        RECT 51.390 41.090 51.740 43.250 ;
        RECT 52.220 41.090 52.570 43.250 ;
        RECT 53.050 41.090 53.400 43.250 ;
        RECT 53.880 41.090 54.230 43.250 ;
        RECT 62.650 42.070 62.820 46.110 ;
        RECT 63.940 42.070 64.110 46.110 ;
        RECT 64.530 42.070 64.700 46.110 ;
        RECT 65.820 42.070 65.990 46.110 ;
        RECT 66.410 42.070 66.580 46.110 ;
        RECT 69.580 42.070 69.750 46.110 ;
        RECT 71.460 42.070 71.630 46.110 ;
        RECT 73.340 42.070 73.510 46.110 ;
        RECT 62.880 41.685 63.880 41.855 ;
        RECT 66.640 41.685 67.640 41.855 ;
        RECT 68.520 41.685 69.520 41.855 ;
        RECT 70.400 41.685 71.400 41.855 ;
        RECT 72.280 41.685 73.280 41.855 ;
        RECT 74.050 41.090 74.400 43.250 ;
        RECT 74.880 41.090 75.230 43.250 ;
        RECT 75.710 41.090 76.060 43.250 ;
        RECT 76.540 41.090 76.890 43.250 ;
        RECT 85.310 42.070 85.480 46.110 ;
        RECT 86.600 42.070 86.770 46.110 ;
        RECT 87.190 42.070 87.360 46.110 ;
        RECT 88.480 42.070 88.650 46.110 ;
        RECT 89.070 42.070 89.240 46.110 ;
        RECT 92.240 42.070 92.410 46.110 ;
        RECT 94.120 42.070 94.290 46.110 ;
        RECT 96.000 42.070 96.170 46.110 ;
        RECT 85.540 41.685 86.540 41.855 ;
        RECT 89.300 41.685 90.300 41.855 ;
        RECT 91.180 41.685 92.180 41.855 ;
        RECT 93.060 41.685 94.060 41.855 ;
        RECT 94.940 41.685 95.940 41.855 ;
        RECT 96.710 41.090 97.060 43.250 ;
        RECT 97.540 41.090 97.890 43.250 ;
        RECT 98.370 41.090 98.720 43.250 ;
        RECT 99.200 41.090 99.550 43.250 ;
        RECT 107.970 42.070 108.140 46.110 ;
        RECT 109.260 42.070 109.430 46.110 ;
        RECT 109.850 42.070 110.020 46.110 ;
        RECT 111.140 42.070 111.310 46.110 ;
        RECT 111.730 42.070 111.900 46.110 ;
        RECT 114.900 42.070 115.070 46.110 ;
        RECT 116.780 42.070 116.950 46.110 ;
        RECT 118.660 42.070 118.830 46.110 ;
        RECT 108.200 41.685 109.200 41.855 ;
        RECT 111.960 41.685 112.960 41.855 ;
        RECT 113.840 41.685 114.840 41.855 ;
        RECT 115.720 41.685 116.720 41.855 ;
        RECT 117.600 41.685 118.600 41.855 ;
        RECT 119.370 41.090 119.720 43.250 ;
        RECT 120.200 41.090 120.550 43.250 ;
        RECT 121.030 41.090 121.380 43.250 ;
        RECT 121.860 41.090 122.210 43.250 ;
      LAYER mcon ;
        RECT 57.565 184.975 57.735 185.145 ;
        RECT 59.405 184.975 59.575 185.145 ;
        RECT 62.625 184.975 62.795 185.145 ;
        RECT 65.845 184.975 66.015 185.145 ;
        RECT 63.545 184.635 63.715 184.805 ;
        RECT 69.525 184.975 69.695 185.145 ;
        RECT 69.985 184.975 70.155 185.145 ;
        RECT 73.205 184.975 73.375 185.145 ;
        RECT 75.965 184.975 76.135 185.145 ;
        RECT 78.265 184.975 78.435 185.145 ;
        RECT 84.245 184.975 84.415 185.145 ;
        RECT 86.545 184.635 86.715 184.805 ;
        RECT 87.465 185.655 87.635 185.825 ;
        RECT 89.305 184.295 89.475 184.465 ;
        RECT 97.125 184.975 97.295 185.145 ;
        RECT 100.805 184.635 100.975 184.805 ;
        RECT 91.145 184.295 91.315 184.465 ;
        RECT 102.185 185.315 102.355 185.485 ;
        RECT 103.105 184.295 103.275 184.465 ;
        RECT 103.565 184.295 103.735 184.465 ;
        RECT 105.405 184.295 105.575 184.465 ;
        RECT 108.165 185.655 108.335 185.825 ;
        RECT 109.545 184.295 109.715 184.465 ;
        RECT 112.305 185.315 112.475 185.485 ;
        RECT 111.845 184.635 112.015 184.805 ;
        RECT 53.425 181.915 53.595 182.085 ;
        RECT 55.265 182.935 55.435 183.105 ;
        RECT 56.645 182.595 56.815 182.765 ;
        RECT 58.025 182.255 58.195 182.425 ;
        RECT 56.185 181.915 56.355 182.085 ;
        RECT 55.265 181.575 55.435 181.745 ;
        RECT 64.465 182.255 64.635 182.425 ;
        RECT 67.225 183.275 67.395 183.445 ;
        RECT 65.385 182.595 65.555 182.765 ;
        RECT 64.925 182.255 65.095 182.425 ;
        RECT 70.445 182.935 70.615 183.105 ;
        RECT 69.525 182.255 69.695 182.425 ;
        RECT 72.745 183.275 72.915 183.445 ;
        RECT 70.905 182.595 71.075 182.765 ;
        RECT 74.585 183.275 74.755 183.445 ;
        RECT 74.125 182.255 74.295 182.425 ;
        RECT 75.045 182.595 75.215 182.765 ;
        RECT 76.885 181.575 77.055 181.745 ;
        RECT 80.105 182.595 80.275 182.765 ;
        RECT 81.485 182.255 81.655 182.425 ;
        RECT 81.945 181.915 82.115 182.085 ;
        RECT 84.245 183.275 84.415 183.445 ;
        RECT 85.165 182.255 85.335 182.425 ;
        RECT 87.925 181.915 88.095 182.085 ;
        RECT 89.765 182.935 89.935 183.105 ;
        RECT 90.225 182.255 90.395 182.425 ;
        RECT 90.685 182.255 90.855 182.425 ;
        RECT 93.905 183.275 94.075 183.445 ;
        RECT 92.065 181.575 92.235 181.745 ;
        RECT 98.045 183.275 98.215 183.445 ;
        RECT 96.205 182.595 96.375 182.765 ;
        RECT 96.665 182.255 96.835 182.425 ;
        RECT 100.345 182.255 100.515 182.425 ;
        RECT 100.805 182.255 100.975 182.425 ;
        RECT 103.105 182.935 103.275 183.105 ;
        RECT 105.865 182.595 106.035 182.765 ;
        RECT 106.785 181.575 106.955 181.745 ;
        RECT 109.085 182.255 109.255 182.425 ;
        RECT 109.545 182.255 109.715 182.425 ;
        RECT 110.925 182.595 111.095 182.765 ;
        RECT 50.665 179.535 50.835 179.705 ;
        RECT 63.085 180.555 63.255 180.725 ;
        RECT 52.045 179.535 52.215 179.705 ;
        RECT 52.965 179.535 53.135 179.705 ;
        RECT 53.885 179.535 54.055 179.705 ;
        RECT 54.345 179.535 54.515 179.705 ;
        RECT 66.305 179.875 66.475 180.045 ;
        RECT 65.385 178.855 65.555 179.025 ;
        RECT 69.065 179.535 69.235 179.705 ;
        RECT 72.745 179.535 72.915 179.705 ;
        RECT 75.965 179.535 76.135 179.705 ;
        RECT 75.045 179.195 75.215 179.365 ;
        RECT 68.145 178.855 68.315 179.025 ;
        RECT 89.765 179.875 89.935 180.045 ;
        RECT 90.225 179.195 90.395 179.365 ;
        RECT 93.905 180.555 94.075 180.725 ;
        RECT 92.985 179.535 93.155 179.705 ;
        RECT 90.685 178.855 90.855 179.025 ;
        RECT 92.525 178.855 92.695 179.025 ;
        RECT 95.745 180.555 95.915 180.725 ;
        RECT 97.125 180.215 97.295 180.385 ;
        RECT 96.665 179.535 96.835 179.705 ;
        RECT 100.345 180.555 100.515 180.725 ;
        RECT 98.505 178.855 98.675 179.025 ;
        RECT 103.105 179.875 103.275 180.045 ;
        RECT 102.645 178.855 102.815 179.025 ;
        RECT 104.485 178.855 104.655 179.025 ;
        RECT 107.245 179.535 107.415 179.705 ;
        RECT 109.085 179.875 109.255 180.045 ;
        RECT 110.465 179.875 110.635 180.045 ;
        RECT 107.705 178.855 107.875 179.025 ;
        RECT 58.485 177.835 58.655 178.005 ;
        RECT 50.665 177.155 50.835 177.325 ;
        RECT 49.745 176.475 49.915 176.645 ;
        RECT 51.585 176.815 51.755 176.985 ;
        RECT 60.785 176.815 60.955 176.985 ;
        RECT 61.245 176.815 61.415 176.985 ;
        RECT 63.545 177.835 63.715 178.005 ;
        RECT 63.085 177.155 63.255 177.325 ;
        RECT 75.965 177.835 76.135 178.005 ;
        RECT 69.065 177.155 69.235 177.325 ;
        RECT 68.145 176.815 68.315 176.985 ;
        RECT 78.265 177.835 78.435 178.005 ;
        RECT 78.725 176.815 78.895 176.985 ;
        RECT 80.105 177.495 80.275 177.665 ;
        RECT 81.480 177.495 81.650 177.665 ;
        RECT 81.895 176.475 82.065 176.645 ;
        RECT 83.325 176.815 83.495 176.985 ;
        RECT 84.120 177.155 84.290 177.325 ;
        RECT 84.705 177.155 84.875 177.325 ;
        RECT 87.000 177.155 87.170 177.325 ;
        RECT 86.085 176.815 86.255 176.985 ;
        RECT 85.125 176.475 85.295 176.645 ;
        RECT 88.385 177.155 88.555 177.325 ;
        RECT 93.905 177.835 94.075 178.005 ;
        RECT 89.765 177.155 89.935 177.325 ;
        RECT 89.305 176.815 89.475 176.985 ;
        RECT 90.685 177.155 90.855 177.325 ;
        RECT 96.205 176.815 96.375 176.985 ;
        RECT 97.125 176.815 97.295 176.985 ;
        RECT 98.505 177.155 98.675 177.325 ;
        RECT 101.265 176.815 101.435 176.985 ;
        RECT 103.105 176.135 103.275 176.305 ;
        RECT 105.405 177.495 105.575 177.665 ;
        RECT 108.165 177.835 108.335 178.005 ;
        RECT 105.865 176.815 106.035 176.985 ;
        RECT 111.385 176.815 111.555 176.985 ;
        RECT 113.685 177.155 113.855 177.325 ;
        RECT 57.565 175.115 57.735 175.285 ;
        RECT 50.205 174.435 50.375 174.605 ;
        RECT 49.745 174.095 49.915 174.265 ;
        RECT 51.585 174.775 51.755 174.945 ;
        RECT 55.725 174.435 55.895 174.605 ;
        RECT 56.185 174.095 56.355 174.265 ;
        RECT 59.405 174.095 59.575 174.265 ;
        RECT 62.625 174.435 62.795 174.605 ;
        RECT 58.485 173.415 58.655 173.585 ;
        RECT 63.545 173.415 63.715 173.585 ;
        RECT 64.005 173.755 64.175 173.925 ;
        RECT 65.845 173.415 66.015 173.585 ;
        RECT 66.305 173.415 66.475 173.585 ;
        RECT 69.065 174.435 69.235 174.605 ;
        RECT 71.135 174.435 71.305 174.605 ;
        RECT 73.665 174.775 73.835 174.945 ;
        RECT 74.625 174.775 74.795 174.945 ;
        RECT 72.750 174.095 72.920 174.265 ;
        RECT 68.605 173.415 68.775 173.585 ;
        RECT 71.830 173.755 72.000 173.925 ;
        RECT 74.590 174.095 74.760 174.265 ;
        RECT 75.630 174.435 75.800 174.605 ;
        RECT 76.425 174.095 76.595 174.265 ;
        RECT 76.935 174.095 77.105 174.265 ;
        RECT 77.855 174.775 78.025 174.945 ;
        RECT 77.350 173.755 77.520 173.925 ;
        RECT 78.775 174.095 78.945 174.265 ;
        RECT 79.645 174.095 79.815 174.265 ;
        RECT 81.945 174.435 82.115 174.605 ;
        RECT 82.405 174.435 82.575 174.605 ;
        RECT 82.865 173.755 83.035 173.925 ;
        RECT 84.705 174.775 84.875 174.945 ;
        RECT 86.085 174.095 86.255 174.265 ;
        RECT 89.305 174.435 89.475 174.605 ;
        RECT 89.765 174.095 89.935 174.265 ;
        RECT 85.165 173.415 85.335 173.585 ;
        RECT 90.225 174.095 90.395 174.265 ;
        RECT 92.065 175.115 92.235 175.285 ;
        RECT 93.445 174.435 93.615 174.605 ;
        RECT 93.905 173.415 94.075 173.585 ;
        RECT 94.365 173.415 94.535 173.585 ;
        RECT 96.205 173.415 96.375 173.585 ;
        RECT 97.585 175.115 97.755 175.285 ;
        RECT 100.805 174.435 100.975 174.605 ;
        RECT 99.885 173.415 100.055 173.585 ;
        RECT 104.025 174.435 104.195 174.605 ;
        RECT 101.725 173.415 101.895 173.585 ;
        RECT 104.485 174.435 104.655 174.605 ;
        RECT 106.785 173.415 106.955 173.585 ;
        RECT 109.545 174.435 109.715 174.605 ;
        RECT 112.765 174.435 112.935 174.605 ;
        RECT 109.085 173.415 109.255 173.585 ;
        RECT 56.185 172.395 56.355 172.565 ;
        RECT 58.485 171.375 58.655 171.545 ;
        RECT 59.405 171.375 59.575 171.545 ;
        RECT 64.005 171.715 64.175 171.885 ;
        RECT 64.925 171.715 65.095 171.885 ;
        RECT 68.145 171.715 68.315 171.885 ;
        RECT 65.845 171.035 66.015 171.205 ;
        RECT 69.065 170.695 69.235 170.865 ;
        RECT 81.025 170.695 81.195 170.865 ;
        RECT 83.325 172.395 83.495 172.565 ;
        RECT 90.225 172.395 90.395 172.565 ;
        RECT 84.245 171.375 84.415 171.545 ;
        RECT 87.005 171.715 87.175 171.885 ;
        RECT 87.925 171.715 88.095 171.885 ;
        RECT 88.385 170.695 88.555 170.865 ;
        RECT 98.045 171.715 98.215 171.885 ;
        RECT 101.725 172.055 101.895 172.225 ;
        RECT 98.965 171.715 99.135 171.885 ;
        RECT 106.330 172.055 106.500 172.225 ;
        RECT 99.425 170.695 99.595 170.865 ;
        RECT 105.865 171.715 106.035 171.885 ;
        RECT 107.250 171.715 107.420 171.885 ;
        RECT 109.545 171.715 109.715 171.885 ;
        RECT 110.130 171.375 110.300 171.545 ;
        RECT 110.925 171.375 111.095 171.545 ;
        RECT 111.850 172.055 112.020 172.225 ;
        RECT 111.435 171.715 111.605 171.885 ;
        RECT 108.165 171.035 108.335 171.205 ;
        RECT 109.125 171.035 109.295 171.205 ;
        RECT 114.145 172.395 114.315 172.565 ;
        RECT 113.275 171.715 113.445 171.885 ;
        RECT 112.355 171.035 112.525 171.205 ;
        RECT 60.785 168.995 60.955 169.165 ;
        RECT 61.705 167.975 61.875 168.145 ;
        RECT 64.005 169.675 64.175 169.845 ;
        RECT 62.165 167.975 62.335 168.145 ;
        RECT 70.905 169.675 71.075 169.845 ;
        RECT 68.145 168.655 68.315 168.825 ;
        RECT 68.605 168.655 68.775 168.825 ;
        RECT 69.525 168.655 69.695 168.825 ;
        RECT 71.825 167.975 71.995 168.145 ;
        RECT 74.585 168.995 74.755 169.165 ;
        RECT 74.125 168.655 74.295 168.825 ;
        RECT 82.865 168.655 83.035 168.825 ;
        RECT 86.125 169.335 86.295 169.505 ;
        RECT 85.165 168.995 85.335 169.165 ;
        RECT 84.250 168.655 84.420 168.825 ;
        RECT 83.330 168.315 83.500 168.485 ;
        RECT 86.090 168.655 86.260 168.825 ;
        RECT 87.130 168.995 87.300 169.165 ;
        RECT 87.925 168.655 88.095 168.825 ;
        RECT 88.435 168.655 88.605 168.825 ;
        RECT 89.355 169.335 89.525 169.505 ;
        RECT 91.145 169.675 91.315 169.845 ;
        RECT 88.850 168.315 89.020 168.485 ;
        RECT 90.275 168.655 90.445 168.825 ;
        RECT 95.745 169.675 95.915 169.845 ;
        RECT 92.985 168.995 93.155 169.165 ;
        RECT 93.445 168.655 93.615 168.825 ;
        RECT 94.365 168.655 94.535 168.825 ;
        RECT 97.585 168.995 97.755 169.165 ;
        RECT 100.845 169.335 101.015 169.505 ;
        RECT 99.885 168.995 100.055 169.165 ;
        RECT 98.970 168.655 99.140 168.825 ;
        RECT 98.050 168.315 98.220 168.485 ;
        RECT 100.810 168.655 100.980 168.825 ;
        RECT 101.850 168.655 102.020 168.825 ;
        RECT 102.645 168.655 102.815 168.825 ;
        RECT 103.155 168.655 103.325 168.825 ;
        RECT 104.075 169.335 104.245 169.505 ;
        RECT 103.570 168.315 103.740 168.485 ;
        RECT 104.995 168.655 105.165 168.825 ;
        RECT 105.865 169.335 106.035 169.505 ;
        RECT 106.785 169.675 106.955 169.845 ;
        RECT 109.545 168.995 109.715 169.165 ;
        RECT 109.085 168.655 109.255 168.825 ;
        RECT 110.925 169.335 111.095 169.505 ;
        RECT 112.305 169.335 112.475 169.505 ;
        RECT 50.665 166.955 50.835 167.125 ;
        RECT 52.040 166.615 52.210 166.785 ;
        RECT 52.455 165.595 52.625 165.765 ;
        RECT 53.885 165.935 54.055 166.105 ;
        RECT 54.680 166.275 54.850 166.445 ;
        RECT 55.265 166.275 55.435 166.445 ;
        RECT 71.365 166.955 71.535 167.125 ;
        RECT 57.560 166.275 57.730 166.445 ;
        RECT 55.685 165.595 55.855 165.765 ;
        RECT 56.645 165.595 56.815 165.765 ;
        RECT 59.175 166.275 59.345 166.445 ;
        RECT 59.865 165.935 60.035 166.105 ;
        RECT 71.825 166.615 71.995 166.785 ;
        RECT 75.965 166.275 76.135 166.445 ;
        RECT 76.885 166.615 77.055 166.785 ;
        RECT 77.805 165.935 77.975 166.105 ;
        RECT 80.565 166.615 80.735 166.785 ;
        RECT 79.645 166.275 79.815 166.445 ;
        RECT 92.525 166.275 92.695 166.445 ;
        RECT 91.605 165.595 91.775 165.765 ;
        RECT 97.125 166.955 97.295 167.125 ;
        RECT 94.825 166.275 94.995 166.445 ;
        RECT 95.745 166.275 95.915 166.445 ;
        RECT 104.945 166.955 105.115 167.125 ;
        RECT 94.365 165.935 94.535 166.105 ;
        RECT 107.245 166.275 107.415 166.445 ;
        RECT 108.165 165.935 108.335 166.105 ;
        RECT 106.785 165.255 106.955 165.425 ;
        RECT 110.005 165.255 110.175 165.425 ;
        RECT 111.845 166.615 112.015 166.785 ;
        RECT 112.305 166.275 112.475 166.445 ;
        RECT 112.765 165.935 112.935 166.105 ;
        RECT 61.245 164.235 61.415 164.405 ;
        RECT 56.645 163.555 56.815 163.725 ;
        RECT 57.105 163.215 57.275 163.385 ;
        RECT 55.265 162.535 55.435 162.705 ;
        RECT 63.035 163.895 63.205 164.065 ;
        RECT 62.620 162.875 62.790 163.045 ;
        RECT 66.265 163.895 66.435 164.065 ;
        RECT 67.225 163.895 67.395 164.065 ;
        RECT 64.465 163.555 64.635 163.725 ;
        RECT 65.260 163.215 65.430 163.385 ;
        RECT 65.845 163.215 66.015 163.385 ;
        RECT 66.300 163.215 66.470 163.385 ;
        RECT 69.525 163.555 69.695 163.725 ;
        RECT 70.445 163.215 70.615 163.385 ;
        RECT 79.645 162.875 79.815 163.045 ;
        RECT 79.185 162.535 79.355 162.705 ;
        RECT 84.245 164.235 84.415 164.405 ;
        RECT 81.485 163.215 81.655 163.385 ;
        RECT 81.945 163.215 82.115 163.385 ;
        RECT 82.865 163.215 83.035 163.385 ;
        RECT 86.085 162.535 86.255 162.705 ;
        RECT 88.845 163.555 89.015 163.725 ;
        RECT 88.385 163.215 88.555 163.385 ;
        RECT 93.905 164.235 94.075 164.405 ;
        RECT 96.665 163.555 96.835 163.725 ;
        RECT 96.205 163.215 96.375 163.385 ;
        RECT 98.045 162.535 98.215 162.705 ;
        RECT 100.805 163.555 100.975 163.725 ;
        RECT 103.105 164.235 103.275 164.405 ;
        RECT 100.345 162.535 100.515 162.705 ;
        RECT 102.645 162.875 102.815 163.045 ;
        RECT 109.545 163.895 109.715 164.065 ;
        RECT 110.465 163.215 110.635 163.385 ;
        RECT 112.305 164.235 112.475 164.405 ;
        RECT 110.925 162.535 111.095 162.705 ;
        RECT 52.965 160.835 53.135 161.005 ;
        RECT 53.425 160.495 53.595 160.665 ;
        RECT 58.025 161.515 58.195 161.685 ;
        RECT 54.805 160.495 54.975 160.665 ;
        RECT 56.185 160.835 56.355 161.005 ;
        RECT 55.725 160.495 55.895 160.665 ;
        RECT 62.165 160.835 62.335 161.005 ;
        RECT 62.625 160.495 62.795 160.665 ;
        RECT 64.005 160.155 64.175 160.325 ;
        RECT 65.385 160.835 65.555 161.005 ;
        RECT 65.845 160.495 66.015 160.665 ;
        RECT 69.985 161.515 70.155 161.685 ;
        RECT 67.225 159.815 67.395 159.985 ;
        RECT 74.125 161.515 74.295 161.685 ;
        RECT 72.285 160.495 72.455 160.665 ;
        RECT 73.205 160.495 73.375 160.665 ;
        RECT 76.425 160.495 76.595 160.665 ;
        RECT 76.885 160.495 77.055 160.665 ;
        RECT 80.105 160.835 80.275 161.005 ;
        RECT 79.645 160.495 79.815 160.665 ;
        RECT 91.605 160.835 91.775 161.005 ;
        RECT 81.485 159.815 81.655 159.985 ;
        RECT 92.065 160.495 92.235 160.665 ;
        RECT 89.765 159.815 89.935 159.985 ;
        RECT 96.665 161.175 96.835 161.345 ;
        RECT 95.745 160.155 95.915 160.325 ;
        RECT 101.725 161.515 101.895 161.685 ;
        RECT 104.025 161.175 104.195 161.345 ;
        RECT 105.865 161.515 106.035 161.685 ;
        RECT 104.485 160.495 104.655 160.665 ;
        RECT 106.785 161.175 106.955 161.345 ;
        RECT 107.705 160.495 107.875 160.665 ;
        RECT 108.625 160.155 108.795 160.325 ;
        RECT 110.925 161.515 111.095 161.685 ;
        RECT 112.305 161.515 112.475 161.685 ;
        RECT 44.685 158.795 44.855 158.965 ;
        RECT 43.765 157.775 43.935 157.945 ;
        RECT 49.745 158.455 49.915 158.625 ;
        RECT 48.825 157.775 48.995 157.945 ;
        RECT 56.185 158.795 56.355 158.965 ;
        RECT 55.265 157.775 55.435 157.945 ;
        RECT 59.865 158.795 60.035 158.965 ;
        RECT 58.945 157.775 59.115 157.945 ;
        RECT 64.925 158.795 65.095 158.965 ;
        RECT 70.445 158.795 70.615 158.965 ;
        RECT 64.005 157.775 64.175 157.945 ;
        RECT 68.605 158.115 68.775 158.285 ;
        RECT 69.065 157.775 69.235 157.945 ;
        RECT 71.365 157.775 71.535 157.945 ;
        RECT 75.045 158.795 75.215 158.965 ;
        RECT 74.125 157.775 74.295 157.945 ;
        RECT 72.285 157.095 72.455 157.265 ;
        RECT 79.185 158.795 79.355 158.965 ;
        RECT 80.105 157.775 80.275 157.945 ;
        RECT 84.705 158.115 84.875 158.285 ;
        RECT 85.165 157.775 85.335 157.945 ;
        RECT 87.465 158.795 87.635 158.965 ;
        RECT 86.545 157.775 86.715 157.945 ;
        RECT 83.325 157.095 83.495 157.265 ;
        RECT 90.225 158.795 90.395 158.965 ;
        RECT 89.305 157.775 89.475 157.945 ;
        RECT 95.285 158.795 95.455 158.965 ;
        RECT 94.365 157.775 94.535 157.945 ;
        RECT 100.345 158.795 100.515 158.965 ;
        RECT 99.425 157.775 99.595 157.945 ;
        RECT 105.405 158.795 105.575 158.965 ;
        RECT 104.485 157.775 104.655 157.945 ;
        RECT 110.005 158.795 110.175 158.965 ;
        RECT 109.545 158.115 109.715 158.285 ;
        RECT 107.705 157.775 107.875 157.945 ;
        RECT 108.625 157.775 108.795 157.945 ;
        RECT 110.925 157.775 111.095 157.945 ;
        RECT 111.845 157.095 112.015 157.265 ;
        RECT 113.225 158.795 113.395 158.965 ;
        RECT 114.145 157.775 114.315 157.945 ;
        RECT 62.960 127.720 63.800 127.890 ;
        RECT 64.840 127.720 65.680 127.890 ;
        RECT 66.720 127.720 67.560 127.890 ;
        RECT 68.600 127.720 69.440 127.890 ;
        RECT 70.480 127.720 71.320 127.890 ;
        RECT 72.360 127.720 73.200 127.890 ;
        RECT 74.240 127.720 75.080 127.890 ;
        RECT 85.620 127.720 86.460 127.890 ;
        RECT 87.500 127.720 88.340 127.890 ;
        RECT 89.380 127.720 90.220 127.890 ;
        RECT 91.260 127.720 92.100 127.890 ;
        RECT 93.140 127.720 93.980 127.890 ;
        RECT 95.020 127.720 95.860 127.890 ;
        RECT 96.900 127.720 97.740 127.890 ;
        RECT 108.280 127.720 109.120 127.890 ;
        RECT 110.160 127.720 111.000 127.890 ;
        RECT 112.040 127.720 112.880 127.890 ;
        RECT 113.920 127.720 114.760 127.890 ;
        RECT 115.800 127.720 116.640 127.890 ;
        RECT 117.680 127.720 118.520 127.890 ;
        RECT 119.560 127.720 120.400 127.890 ;
        RECT 62.650 125.590 62.820 127.470 ;
        RECT 65.820 125.590 65.990 127.470 ;
        RECT 66.410 125.590 66.580 127.470 ;
        RECT 67.700 125.590 67.870 127.470 ;
        RECT 68.290 125.590 68.460 127.470 ;
        RECT 69.580 125.590 69.750 127.470 ;
        RECT 71.460 125.590 71.630 127.470 ;
        RECT 73.340 125.590 73.510 127.470 ;
        RECT 75.220 125.590 75.390 127.470 ;
        RECT 62.960 125.170 63.800 125.340 ;
        RECT 64.840 125.170 65.680 125.340 ;
        RECT 66.720 125.170 67.560 125.340 ;
        RECT 68.600 125.170 69.440 125.340 ;
        RECT 70.480 125.170 71.320 125.340 ;
        RECT 72.360 125.170 73.200 125.340 ;
        RECT 74.240 125.170 75.080 125.340 ;
        RECT 62.960 124.630 63.800 124.800 ;
        RECT 64.840 124.630 65.680 124.800 ;
        RECT 66.720 124.630 67.560 124.800 ;
        RECT 68.600 124.630 69.440 124.800 ;
        RECT 70.480 124.630 71.320 124.800 ;
        RECT 72.360 124.630 73.200 124.800 ;
        RECT 74.240 124.630 75.080 124.800 ;
        RECT 62.650 122.500 62.820 124.380 ;
        RECT 58.990 122.330 59.330 122.500 ;
        RECT 60.390 122.330 60.730 122.500 ;
        RECT 65.820 122.500 65.990 124.380 ;
        RECT 66.410 122.500 66.580 124.380 ;
        RECT 67.700 122.500 67.870 124.380 ;
        RECT 68.290 122.500 68.460 124.380 ;
        RECT 69.580 122.500 69.750 124.380 ;
        RECT 71.460 122.500 71.630 124.380 ;
        RECT 73.340 122.500 73.510 124.380 ;
        RECT 75.220 122.500 75.390 124.380 ;
        RECT 58.680 121.700 58.850 122.080 ;
        RECT 62.960 122.080 63.800 122.250 ;
        RECT 64.840 122.080 65.680 122.250 ;
        RECT 66.720 122.080 67.560 122.250 ;
        RECT 68.600 122.080 69.440 122.250 ;
        RECT 70.480 122.080 71.320 122.250 ;
        RECT 72.360 122.080 73.200 122.250 ;
        RECT 74.240 122.080 75.080 122.250 ;
        RECT 60.080 121.700 60.250 122.080 ;
        RECT 62.960 121.525 63.800 121.695 ;
        RECT 64.840 121.525 65.680 121.695 ;
        RECT 66.720 121.525 67.560 121.695 ;
        RECT 68.600 121.525 69.440 121.695 ;
        RECT 70.480 121.525 71.320 121.695 ;
        RECT 72.360 121.525 73.200 121.695 ;
        RECT 58.990 121.280 59.330 121.450 ;
        RECT 60.390 121.280 60.730 121.450 ;
        RECT 58.990 120.715 59.330 120.885 ;
        RECT 60.390 120.715 60.730 120.885 ;
        RECT 58.680 119.540 58.850 120.420 ;
        RECT 60.080 119.540 60.250 120.420 ;
        RECT 58.990 119.075 59.330 119.245 ;
        RECT 60.390 119.075 60.730 119.245 ;
        RECT 62.650 117.350 62.820 121.230 ;
        RECT 63.940 117.350 64.110 121.230 ;
        RECT 64.530 117.350 64.700 121.230 ;
        RECT 65.820 117.350 65.990 121.230 ;
        RECT 66.410 117.350 66.580 121.230 ;
        RECT 69.580 117.350 69.750 121.230 ;
        RECT 71.460 117.350 71.630 121.230 ;
        RECT 73.340 117.350 73.510 121.230 ;
        RECT 74.130 119.445 74.320 121.430 ;
        RECT 74.960 119.445 75.150 121.430 ;
        RECT 75.790 119.445 75.980 121.430 ;
        RECT 78.960 124.705 79.150 126.690 ;
        RECT 78.960 120.210 79.150 122.195 ;
        RECT 85.310 125.590 85.480 127.470 ;
        RECT 88.480 125.590 88.650 127.470 ;
        RECT 89.070 125.590 89.240 127.470 ;
        RECT 90.360 125.590 90.530 127.470 ;
        RECT 90.950 125.590 91.120 127.470 ;
        RECT 92.240 125.590 92.410 127.470 ;
        RECT 94.120 125.590 94.290 127.470 ;
        RECT 96.000 125.590 96.170 127.470 ;
        RECT 97.880 125.590 98.050 127.470 ;
        RECT 85.620 125.170 86.460 125.340 ;
        RECT 87.500 125.170 88.340 125.340 ;
        RECT 89.380 125.170 90.220 125.340 ;
        RECT 91.260 125.170 92.100 125.340 ;
        RECT 93.140 125.170 93.980 125.340 ;
        RECT 95.020 125.170 95.860 125.340 ;
        RECT 96.900 125.170 97.740 125.340 ;
        RECT 85.620 124.630 86.460 124.800 ;
        RECT 87.500 124.630 88.340 124.800 ;
        RECT 89.380 124.630 90.220 124.800 ;
        RECT 91.260 124.630 92.100 124.800 ;
        RECT 93.140 124.630 93.980 124.800 ;
        RECT 95.020 124.630 95.860 124.800 ;
        RECT 96.900 124.630 97.740 124.800 ;
        RECT 85.310 122.500 85.480 124.380 ;
        RECT 81.650 122.330 81.990 122.500 ;
        RECT 83.050 122.330 83.390 122.500 ;
        RECT 88.480 122.500 88.650 124.380 ;
        RECT 89.070 122.500 89.240 124.380 ;
        RECT 90.360 122.500 90.530 124.380 ;
        RECT 90.950 122.500 91.120 124.380 ;
        RECT 92.240 122.500 92.410 124.380 ;
        RECT 94.120 122.500 94.290 124.380 ;
        RECT 96.000 122.500 96.170 124.380 ;
        RECT 97.880 122.500 98.050 124.380 ;
        RECT 81.340 121.700 81.510 122.080 ;
        RECT 85.620 122.080 86.460 122.250 ;
        RECT 87.500 122.080 88.340 122.250 ;
        RECT 89.380 122.080 90.220 122.250 ;
        RECT 91.260 122.080 92.100 122.250 ;
        RECT 93.140 122.080 93.980 122.250 ;
        RECT 95.020 122.080 95.860 122.250 ;
        RECT 96.900 122.080 97.740 122.250 ;
        RECT 82.740 121.700 82.910 122.080 ;
        RECT 85.620 121.525 86.460 121.695 ;
        RECT 87.500 121.525 88.340 121.695 ;
        RECT 89.380 121.525 90.220 121.695 ;
        RECT 91.260 121.525 92.100 121.695 ;
        RECT 93.140 121.525 93.980 121.695 ;
        RECT 95.020 121.525 95.860 121.695 ;
        RECT 81.650 121.280 81.990 121.450 ;
        RECT 83.050 121.280 83.390 121.450 ;
        RECT 81.650 120.715 81.990 120.885 ;
        RECT 83.050 120.715 83.390 120.885 ;
        RECT 62.960 116.885 63.800 117.055 ;
        RECT 64.840 116.885 65.680 117.055 ;
        RECT 66.720 116.885 67.560 117.055 ;
        RECT 68.600 116.885 69.440 117.055 ;
        RECT 70.480 116.885 71.320 117.055 ;
        RECT 72.360 116.885 73.200 117.055 ;
        RECT 62.960 116.345 63.800 116.515 ;
        RECT 64.840 116.345 65.680 116.515 ;
        RECT 66.720 116.345 67.560 116.515 ;
        RECT 68.600 116.345 69.440 116.515 ;
        RECT 70.480 116.345 71.320 116.515 ;
        RECT 72.360 116.345 73.200 116.515 ;
        RECT 62.650 112.170 62.820 116.050 ;
        RECT 63.940 112.170 64.110 116.050 ;
        RECT 64.530 112.170 64.700 116.050 ;
        RECT 65.820 112.170 65.990 116.050 ;
        RECT 66.410 112.170 66.580 116.050 ;
        RECT 69.580 112.170 69.750 116.050 ;
        RECT 71.460 112.170 71.630 116.050 ;
        RECT 73.340 112.170 73.510 116.050 ;
        RECT 62.960 111.705 63.800 111.875 ;
        RECT 64.840 111.705 65.680 111.875 ;
        RECT 66.720 111.705 67.560 111.875 ;
        RECT 68.600 111.705 69.440 111.875 ;
        RECT 70.480 111.705 71.320 111.875 ;
        RECT 72.360 111.705 73.200 111.875 ;
        RECT 74.130 111.200 74.320 113.185 ;
        RECT 74.960 111.200 75.150 113.185 ;
        RECT 75.790 111.200 75.980 113.185 ;
        RECT 76.620 111.200 76.810 113.185 ;
        RECT 78.960 116.915 79.150 118.900 ;
        RECT 78.960 112.420 79.150 114.405 ;
        RECT 81.340 119.540 81.510 120.420 ;
        RECT 82.740 119.540 82.910 120.420 ;
        RECT 81.650 119.075 81.990 119.245 ;
        RECT 83.050 119.075 83.390 119.245 ;
        RECT 85.310 117.350 85.480 121.230 ;
        RECT 86.600 117.350 86.770 121.230 ;
        RECT 87.190 117.350 87.360 121.230 ;
        RECT 88.480 117.350 88.650 121.230 ;
        RECT 89.070 117.350 89.240 121.230 ;
        RECT 92.240 117.350 92.410 121.230 ;
        RECT 94.120 117.350 94.290 121.230 ;
        RECT 96.000 117.350 96.170 121.230 ;
        RECT 96.790 119.445 96.980 121.430 ;
        RECT 97.620 119.445 97.810 121.430 ;
        RECT 98.450 119.445 98.640 121.430 ;
        RECT 101.620 124.705 101.810 126.690 ;
        RECT 101.620 120.210 101.810 122.195 ;
        RECT 107.970 125.590 108.140 127.470 ;
        RECT 111.140 125.590 111.310 127.470 ;
        RECT 111.730 125.590 111.900 127.470 ;
        RECT 113.020 125.590 113.190 127.470 ;
        RECT 113.610 125.590 113.780 127.470 ;
        RECT 114.900 125.590 115.070 127.470 ;
        RECT 116.780 125.590 116.950 127.470 ;
        RECT 118.660 125.590 118.830 127.470 ;
        RECT 120.540 125.590 120.710 127.470 ;
        RECT 108.280 125.170 109.120 125.340 ;
        RECT 110.160 125.170 111.000 125.340 ;
        RECT 112.040 125.170 112.880 125.340 ;
        RECT 113.920 125.170 114.760 125.340 ;
        RECT 115.800 125.170 116.640 125.340 ;
        RECT 117.680 125.170 118.520 125.340 ;
        RECT 119.560 125.170 120.400 125.340 ;
        RECT 108.280 124.630 109.120 124.800 ;
        RECT 110.160 124.630 111.000 124.800 ;
        RECT 112.040 124.630 112.880 124.800 ;
        RECT 113.920 124.630 114.760 124.800 ;
        RECT 115.800 124.630 116.640 124.800 ;
        RECT 117.680 124.630 118.520 124.800 ;
        RECT 119.560 124.630 120.400 124.800 ;
        RECT 107.970 122.500 108.140 124.380 ;
        RECT 104.310 122.330 104.650 122.500 ;
        RECT 105.710 122.330 106.050 122.500 ;
        RECT 111.140 122.500 111.310 124.380 ;
        RECT 111.730 122.500 111.900 124.380 ;
        RECT 113.020 122.500 113.190 124.380 ;
        RECT 113.610 122.500 113.780 124.380 ;
        RECT 114.900 122.500 115.070 124.380 ;
        RECT 116.780 122.500 116.950 124.380 ;
        RECT 118.660 122.500 118.830 124.380 ;
        RECT 120.540 122.500 120.710 124.380 ;
        RECT 104.000 121.700 104.170 122.080 ;
        RECT 108.280 122.080 109.120 122.250 ;
        RECT 110.160 122.080 111.000 122.250 ;
        RECT 112.040 122.080 112.880 122.250 ;
        RECT 113.920 122.080 114.760 122.250 ;
        RECT 115.800 122.080 116.640 122.250 ;
        RECT 117.680 122.080 118.520 122.250 ;
        RECT 119.560 122.080 120.400 122.250 ;
        RECT 105.400 121.700 105.570 122.080 ;
        RECT 108.280 121.525 109.120 121.695 ;
        RECT 110.160 121.525 111.000 121.695 ;
        RECT 112.040 121.525 112.880 121.695 ;
        RECT 113.920 121.525 114.760 121.695 ;
        RECT 115.800 121.525 116.640 121.695 ;
        RECT 117.680 121.525 118.520 121.695 ;
        RECT 104.310 121.280 104.650 121.450 ;
        RECT 105.710 121.280 106.050 121.450 ;
        RECT 104.310 120.715 104.650 120.885 ;
        RECT 105.710 120.715 106.050 120.885 ;
        RECT 85.620 116.885 86.460 117.055 ;
        RECT 87.500 116.885 88.340 117.055 ;
        RECT 89.380 116.885 90.220 117.055 ;
        RECT 91.260 116.885 92.100 117.055 ;
        RECT 93.140 116.885 93.980 117.055 ;
        RECT 95.020 116.885 95.860 117.055 ;
        RECT 85.620 116.345 86.460 116.515 ;
        RECT 87.500 116.345 88.340 116.515 ;
        RECT 89.380 116.345 90.220 116.515 ;
        RECT 91.260 116.345 92.100 116.515 ;
        RECT 93.140 116.345 93.980 116.515 ;
        RECT 95.020 116.345 95.860 116.515 ;
        RECT 85.310 112.170 85.480 116.050 ;
        RECT 86.600 112.170 86.770 116.050 ;
        RECT 87.190 112.170 87.360 116.050 ;
        RECT 88.480 112.170 88.650 116.050 ;
        RECT 89.070 112.170 89.240 116.050 ;
        RECT 92.240 112.170 92.410 116.050 ;
        RECT 94.120 112.170 94.290 116.050 ;
        RECT 96.000 112.170 96.170 116.050 ;
        RECT 85.620 111.705 86.460 111.875 ;
        RECT 87.500 111.705 88.340 111.875 ;
        RECT 89.380 111.705 90.220 111.875 ;
        RECT 91.260 111.705 92.100 111.875 ;
        RECT 93.140 111.705 93.980 111.875 ;
        RECT 95.020 111.705 95.860 111.875 ;
        RECT 96.790 111.200 96.980 113.185 ;
        RECT 97.620 111.200 97.810 113.185 ;
        RECT 98.450 111.200 98.640 113.185 ;
        RECT 99.280 111.200 99.470 113.185 ;
        RECT 101.620 116.915 101.810 118.900 ;
        RECT 101.620 112.420 101.810 114.405 ;
        RECT 104.000 119.540 104.170 120.420 ;
        RECT 105.400 119.540 105.570 120.420 ;
        RECT 104.310 119.075 104.650 119.245 ;
        RECT 105.710 119.075 106.050 119.245 ;
        RECT 107.970 117.350 108.140 121.230 ;
        RECT 109.260 117.350 109.430 121.230 ;
        RECT 109.850 117.350 110.020 121.230 ;
        RECT 111.140 117.350 111.310 121.230 ;
        RECT 111.730 117.350 111.900 121.230 ;
        RECT 114.900 117.350 115.070 121.230 ;
        RECT 116.780 117.350 116.950 121.230 ;
        RECT 118.660 117.350 118.830 121.230 ;
        RECT 119.450 119.445 119.640 121.430 ;
        RECT 120.280 119.445 120.470 121.430 ;
        RECT 121.110 119.445 121.300 121.430 ;
        RECT 124.280 120.210 124.470 122.195 ;
        RECT 108.280 116.885 109.120 117.055 ;
        RECT 110.160 116.885 111.000 117.055 ;
        RECT 112.040 116.885 112.880 117.055 ;
        RECT 113.920 116.885 114.760 117.055 ;
        RECT 115.800 116.885 116.640 117.055 ;
        RECT 117.680 116.885 118.520 117.055 ;
        RECT 108.280 116.345 109.120 116.515 ;
        RECT 110.160 116.345 111.000 116.515 ;
        RECT 112.040 116.345 112.880 116.515 ;
        RECT 113.920 116.345 114.760 116.515 ;
        RECT 115.800 116.345 116.640 116.515 ;
        RECT 117.680 116.345 118.520 116.515 ;
        RECT 107.970 112.170 108.140 116.050 ;
        RECT 109.260 112.170 109.430 116.050 ;
        RECT 109.850 112.170 110.020 116.050 ;
        RECT 111.140 112.170 111.310 116.050 ;
        RECT 111.730 112.170 111.900 116.050 ;
        RECT 114.900 112.170 115.070 116.050 ;
        RECT 116.780 112.170 116.950 116.050 ;
        RECT 118.660 112.170 118.830 116.050 ;
        RECT 108.280 111.705 109.120 111.875 ;
        RECT 110.160 111.705 111.000 111.875 ;
        RECT 112.040 111.705 112.880 111.875 ;
        RECT 113.920 111.705 114.760 111.875 ;
        RECT 115.800 111.705 116.640 111.875 ;
        RECT 117.680 111.705 118.520 111.875 ;
        RECT 119.450 111.200 119.640 113.185 ;
        RECT 120.280 111.200 120.470 113.185 ;
        RECT 121.110 111.200 121.300 113.185 ;
        RECT 121.940 111.200 122.130 113.185 ;
        RECT 124.280 116.915 124.470 118.900 ;
        RECT 124.280 112.420 124.470 114.405 ;
        RECT 40.300 110.380 41.140 110.550 ;
        RECT 42.180 110.380 43.020 110.550 ;
        RECT 44.060 110.380 44.900 110.550 ;
        RECT 45.940 110.380 46.780 110.550 ;
        RECT 47.820 110.380 48.660 110.550 ;
        RECT 49.700 110.380 50.540 110.550 ;
        RECT 51.580 110.380 52.420 110.550 ;
        RECT 62.960 110.380 63.800 110.550 ;
        RECT 64.840 110.380 65.680 110.550 ;
        RECT 66.720 110.380 67.560 110.550 ;
        RECT 68.600 110.380 69.440 110.550 ;
        RECT 70.480 110.380 71.320 110.550 ;
        RECT 72.360 110.380 73.200 110.550 ;
        RECT 74.240 110.380 75.080 110.550 ;
        RECT 85.620 110.380 86.460 110.550 ;
        RECT 87.500 110.380 88.340 110.550 ;
        RECT 89.380 110.380 90.220 110.550 ;
        RECT 91.260 110.380 92.100 110.550 ;
        RECT 93.140 110.380 93.980 110.550 ;
        RECT 95.020 110.380 95.860 110.550 ;
        RECT 96.900 110.380 97.740 110.550 ;
        RECT 108.280 110.380 109.120 110.550 ;
        RECT 110.160 110.380 111.000 110.550 ;
        RECT 112.040 110.380 112.880 110.550 ;
        RECT 113.920 110.380 114.760 110.550 ;
        RECT 115.800 110.380 116.640 110.550 ;
        RECT 117.680 110.380 118.520 110.550 ;
        RECT 119.560 110.380 120.400 110.550 ;
        RECT 39.990 108.250 40.160 110.130 ;
        RECT 43.160 108.250 43.330 110.130 ;
        RECT 43.750 108.250 43.920 110.130 ;
        RECT 45.040 108.250 45.210 110.130 ;
        RECT 45.630 108.250 45.800 110.130 ;
        RECT 46.920 108.250 47.090 110.130 ;
        RECT 48.800 108.250 48.970 110.130 ;
        RECT 50.680 108.250 50.850 110.130 ;
        RECT 52.560 108.250 52.730 110.130 ;
        RECT 40.300 107.830 41.140 108.000 ;
        RECT 42.180 107.830 43.020 108.000 ;
        RECT 44.060 107.830 44.900 108.000 ;
        RECT 45.940 107.830 46.780 108.000 ;
        RECT 47.820 107.830 48.660 108.000 ;
        RECT 49.700 107.830 50.540 108.000 ;
        RECT 51.580 107.830 52.420 108.000 ;
        RECT 40.300 107.290 41.140 107.460 ;
        RECT 42.180 107.290 43.020 107.460 ;
        RECT 44.060 107.290 44.900 107.460 ;
        RECT 45.940 107.290 46.780 107.460 ;
        RECT 47.820 107.290 48.660 107.460 ;
        RECT 49.700 107.290 50.540 107.460 ;
        RECT 51.580 107.290 52.420 107.460 ;
        RECT 39.990 105.160 40.160 107.040 ;
        RECT 36.330 104.990 36.670 105.160 ;
        RECT 37.730 104.990 38.070 105.160 ;
        RECT 43.160 105.160 43.330 107.040 ;
        RECT 43.750 105.160 43.920 107.040 ;
        RECT 45.040 105.160 45.210 107.040 ;
        RECT 45.630 105.160 45.800 107.040 ;
        RECT 46.920 105.160 47.090 107.040 ;
        RECT 48.800 105.160 48.970 107.040 ;
        RECT 50.680 105.160 50.850 107.040 ;
        RECT 52.560 105.160 52.730 107.040 ;
        RECT 36.020 104.360 36.190 104.740 ;
        RECT 40.300 104.740 41.140 104.910 ;
        RECT 42.180 104.740 43.020 104.910 ;
        RECT 44.060 104.740 44.900 104.910 ;
        RECT 45.940 104.740 46.780 104.910 ;
        RECT 47.820 104.740 48.660 104.910 ;
        RECT 49.700 104.740 50.540 104.910 ;
        RECT 51.580 104.740 52.420 104.910 ;
        RECT 37.420 104.360 37.590 104.740 ;
        RECT 40.300 104.185 41.140 104.355 ;
        RECT 42.180 104.185 43.020 104.355 ;
        RECT 44.060 104.185 44.900 104.355 ;
        RECT 45.940 104.185 46.780 104.355 ;
        RECT 47.820 104.185 48.660 104.355 ;
        RECT 49.700 104.185 50.540 104.355 ;
        RECT 36.330 103.940 36.670 104.110 ;
        RECT 37.730 103.940 38.070 104.110 ;
        RECT 36.330 103.375 36.670 103.545 ;
        RECT 37.730 103.375 38.070 103.545 ;
        RECT 36.020 102.200 36.190 103.080 ;
        RECT 37.420 102.200 37.590 103.080 ;
        RECT 36.330 101.735 36.670 101.905 ;
        RECT 37.730 101.735 38.070 101.905 ;
        RECT 39.990 100.010 40.160 103.890 ;
        RECT 41.280 100.010 41.450 103.890 ;
        RECT 41.870 100.010 42.040 103.890 ;
        RECT 43.160 100.010 43.330 103.890 ;
        RECT 43.750 100.010 43.920 103.890 ;
        RECT 46.920 100.010 47.090 103.890 ;
        RECT 48.800 100.010 48.970 103.890 ;
        RECT 50.680 100.010 50.850 103.890 ;
        RECT 51.470 102.105 51.660 104.090 ;
        RECT 52.300 102.105 52.490 104.090 ;
        RECT 53.130 102.105 53.320 104.090 ;
        RECT 56.300 102.870 56.490 104.855 ;
        RECT 62.650 108.250 62.820 110.130 ;
        RECT 65.820 108.250 65.990 110.130 ;
        RECT 66.410 108.250 66.580 110.130 ;
        RECT 67.700 108.250 67.870 110.130 ;
        RECT 68.290 108.250 68.460 110.130 ;
        RECT 69.580 108.250 69.750 110.130 ;
        RECT 71.460 108.250 71.630 110.130 ;
        RECT 73.340 108.250 73.510 110.130 ;
        RECT 75.220 108.250 75.390 110.130 ;
        RECT 62.960 107.830 63.800 108.000 ;
        RECT 64.840 107.830 65.680 108.000 ;
        RECT 66.720 107.830 67.560 108.000 ;
        RECT 68.600 107.830 69.440 108.000 ;
        RECT 70.480 107.830 71.320 108.000 ;
        RECT 72.360 107.830 73.200 108.000 ;
        RECT 74.240 107.830 75.080 108.000 ;
        RECT 62.960 107.290 63.800 107.460 ;
        RECT 64.840 107.290 65.680 107.460 ;
        RECT 66.720 107.290 67.560 107.460 ;
        RECT 68.600 107.290 69.440 107.460 ;
        RECT 70.480 107.290 71.320 107.460 ;
        RECT 72.360 107.290 73.200 107.460 ;
        RECT 74.240 107.290 75.080 107.460 ;
        RECT 62.650 105.160 62.820 107.040 ;
        RECT 58.990 104.990 59.330 105.160 ;
        RECT 60.390 104.990 60.730 105.160 ;
        RECT 65.820 105.160 65.990 107.040 ;
        RECT 66.410 105.160 66.580 107.040 ;
        RECT 67.700 105.160 67.870 107.040 ;
        RECT 68.290 105.160 68.460 107.040 ;
        RECT 69.580 105.160 69.750 107.040 ;
        RECT 71.460 105.160 71.630 107.040 ;
        RECT 73.340 105.160 73.510 107.040 ;
        RECT 75.220 105.160 75.390 107.040 ;
        RECT 58.680 104.360 58.850 104.740 ;
        RECT 62.960 104.740 63.800 104.910 ;
        RECT 64.840 104.740 65.680 104.910 ;
        RECT 66.720 104.740 67.560 104.910 ;
        RECT 68.600 104.740 69.440 104.910 ;
        RECT 70.480 104.740 71.320 104.910 ;
        RECT 72.360 104.740 73.200 104.910 ;
        RECT 74.240 104.740 75.080 104.910 ;
        RECT 60.080 104.360 60.250 104.740 ;
        RECT 62.960 104.185 63.800 104.355 ;
        RECT 64.840 104.185 65.680 104.355 ;
        RECT 66.720 104.185 67.560 104.355 ;
        RECT 68.600 104.185 69.440 104.355 ;
        RECT 70.480 104.185 71.320 104.355 ;
        RECT 72.360 104.185 73.200 104.355 ;
        RECT 58.990 103.940 59.330 104.110 ;
        RECT 60.390 103.940 60.730 104.110 ;
        RECT 58.990 103.375 59.330 103.545 ;
        RECT 60.390 103.375 60.730 103.545 ;
        RECT 40.300 99.545 41.140 99.715 ;
        RECT 42.180 99.545 43.020 99.715 ;
        RECT 44.060 99.545 44.900 99.715 ;
        RECT 45.940 99.545 46.780 99.715 ;
        RECT 47.820 99.545 48.660 99.715 ;
        RECT 49.700 99.545 50.540 99.715 ;
        RECT 40.300 99.005 41.140 99.175 ;
        RECT 42.180 99.005 43.020 99.175 ;
        RECT 44.060 99.005 44.900 99.175 ;
        RECT 45.940 99.005 46.780 99.175 ;
        RECT 47.820 99.005 48.660 99.175 ;
        RECT 49.700 99.005 50.540 99.175 ;
        RECT 39.990 94.830 40.160 98.710 ;
        RECT 41.280 94.830 41.450 98.710 ;
        RECT 41.870 94.830 42.040 98.710 ;
        RECT 43.160 94.830 43.330 98.710 ;
        RECT 43.750 94.830 43.920 98.710 ;
        RECT 46.920 94.830 47.090 98.710 ;
        RECT 48.800 94.830 48.970 98.710 ;
        RECT 50.680 94.830 50.850 98.710 ;
        RECT 40.300 94.365 41.140 94.535 ;
        RECT 42.180 94.365 43.020 94.535 ;
        RECT 44.060 94.365 44.900 94.535 ;
        RECT 45.940 94.365 46.780 94.535 ;
        RECT 47.820 94.365 48.660 94.535 ;
        RECT 49.700 94.365 50.540 94.535 ;
        RECT 51.470 93.860 51.660 95.845 ;
        RECT 52.300 93.860 52.490 95.845 ;
        RECT 53.130 93.860 53.320 95.845 ;
        RECT 53.960 93.860 54.150 95.845 ;
        RECT 56.300 99.575 56.490 101.560 ;
        RECT 56.300 95.080 56.490 97.065 ;
        RECT 58.680 102.200 58.850 103.080 ;
        RECT 60.080 102.200 60.250 103.080 ;
        RECT 58.990 101.735 59.330 101.905 ;
        RECT 60.390 101.735 60.730 101.905 ;
        RECT 62.650 100.010 62.820 103.890 ;
        RECT 63.940 100.010 64.110 103.890 ;
        RECT 64.530 100.010 64.700 103.890 ;
        RECT 65.820 100.010 65.990 103.890 ;
        RECT 66.410 100.010 66.580 103.890 ;
        RECT 69.580 100.010 69.750 103.890 ;
        RECT 71.460 100.010 71.630 103.890 ;
        RECT 73.340 100.010 73.510 103.890 ;
        RECT 74.130 102.105 74.320 104.090 ;
        RECT 74.960 102.105 75.150 104.090 ;
        RECT 75.790 102.105 75.980 104.090 ;
        RECT 78.960 107.365 79.150 109.350 ;
        RECT 78.960 102.870 79.150 104.855 ;
        RECT 85.310 108.250 85.480 110.130 ;
        RECT 88.480 108.250 88.650 110.130 ;
        RECT 89.070 108.250 89.240 110.130 ;
        RECT 90.360 108.250 90.530 110.130 ;
        RECT 90.950 108.250 91.120 110.130 ;
        RECT 92.240 108.250 92.410 110.130 ;
        RECT 94.120 108.250 94.290 110.130 ;
        RECT 96.000 108.250 96.170 110.130 ;
        RECT 97.880 108.250 98.050 110.130 ;
        RECT 85.620 107.830 86.460 108.000 ;
        RECT 87.500 107.830 88.340 108.000 ;
        RECT 89.380 107.830 90.220 108.000 ;
        RECT 91.260 107.830 92.100 108.000 ;
        RECT 93.140 107.830 93.980 108.000 ;
        RECT 95.020 107.830 95.860 108.000 ;
        RECT 96.900 107.830 97.740 108.000 ;
        RECT 85.620 107.290 86.460 107.460 ;
        RECT 87.500 107.290 88.340 107.460 ;
        RECT 89.380 107.290 90.220 107.460 ;
        RECT 91.260 107.290 92.100 107.460 ;
        RECT 93.140 107.290 93.980 107.460 ;
        RECT 95.020 107.290 95.860 107.460 ;
        RECT 96.900 107.290 97.740 107.460 ;
        RECT 85.310 105.160 85.480 107.040 ;
        RECT 81.650 104.990 81.990 105.160 ;
        RECT 83.050 104.990 83.390 105.160 ;
        RECT 88.480 105.160 88.650 107.040 ;
        RECT 89.070 105.160 89.240 107.040 ;
        RECT 90.360 105.160 90.530 107.040 ;
        RECT 90.950 105.160 91.120 107.040 ;
        RECT 92.240 105.160 92.410 107.040 ;
        RECT 94.120 105.160 94.290 107.040 ;
        RECT 96.000 105.160 96.170 107.040 ;
        RECT 97.880 105.160 98.050 107.040 ;
        RECT 81.340 104.360 81.510 104.740 ;
        RECT 85.620 104.740 86.460 104.910 ;
        RECT 87.500 104.740 88.340 104.910 ;
        RECT 89.380 104.740 90.220 104.910 ;
        RECT 91.260 104.740 92.100 104.910 ;
        RECT 93.140 104.740 93.980 104.910 ;
        RECT 95.020 104.740 95.860 104.910 ;
        RECT 96.900 104.740 97.740 104.910 ;
        RECT 82.740 104.360 82.910 104.740 ;
        RECT 85.620 104.185 86.460 104.355 ;
        RECT 87.500 104.185 88.340 104.355 ;
        RECT 89.380 104.185 90.220 104.355 ;
        RECT 91.260 104.185 92.100 104.355 ;
        RECT 93.140 104.185 93.980 104.355 ;
        RECT 95.020 104.185 95.860 104.355 ;
        RECT 81.650 103.940 81.990 104.110 ;
        RECT 83.050 103.940 83.390 104.110 ;
        RECT 81.650 103.375 81.990 103.545 ;
        RECT 83.050 103.375 83.390 103.545 ;
        RECT 62.960 99.545 63.800 99.715 ;
        RECT 64.840 99.545 65.680 99.715 ;
        RECT 66.720 99.545 67.560 99.715 ;
        RECT 68.600 99.545 69.440 99.715 ;
        RECT 70.480 99.545 71.320 99.715 ;
        RECT 72.360 99.545 73.200 99.715 ;
        RECT 62.960 99.005 63.800 99.175 ;
        RECT 64.840 99.005 65.680 99.175 ;
        RECT 66.720 99.005 67.560 99.175 ;
        RECT 68.600 99.005 69.440 99.175 ;
        RECT 70.480 99.005 71.320 99.175 ;
        RECT 72.360 99.005 73.200 99.175 ;
        RECT 62.650 94.830 62.820 98.710 ;
        RECT 63.940 94.830 64.110 98.710 ;
        RECT 64.530 94.830 64.700 98.710 ;
        RECT 65.820 94.830 65.990 98.710 ;
        RECT 66.410 94.830 66.580 98.710 ;
        RECT 69.580 94.830 69.750 98.710 ;
        RECT 71.460 94.830 71.630 98.710 ;
        RECT 73.340 94.830 73.510 98.710 ;
        RECT 62.960 94.365 63.800 94.535 ;
        RECT 64.840 94.365 65.680 94.535 ;
        RECT 66.720 94.365 67.560 94.535 ;
        RECT 68.600 94.365 69.440 94.535 ;
        RECT 70.480 94.365 71.320 94.535 ;
        RECT 72.360 94.365 73.200 94.535 ;
        RECT 74.130 93.860 74.320 95.845 ;
        RECT 74.960 93.860 75.150 95.845 ;
        RECT 75.790 93.860 75.980 95.845 ;
        RECT 76.620 93.860 76.810 95.845 ;
        RECT 78.960 99.575 79.150 101.560 ;
        RECT 78.960 95.080 79.150 97.065 ;
        RECT 81.340 102.200 81.510 103.080 ;
        RECT 82.740 102.200 82.910 103.080 ;
        RECT 81.650 101.735 81.990 101.905 ;
        RECT 83.050 101.735 83.390 101.905 ;
        RECT 85.310 100.010 85.480 103.890 ;
        RECT 86.600 100.010 86.770 103.890 ;
        RECT 87.190 100.010 87.360 103.890 ;
        RECT 88.480 100.010 88.650 103.890 ;
        RECT 89.070 100.010 89.240 103.890 ;
        RECT 92.240 100.010 92.410 103.890 ;
        RECT 94.120 100.010 94.290 103.890 ;
        RECT 96.000 100.010 96.170 103.890 ;
        RECT 96.790 102.105 96.980 104.090 ;
        RECT 97.620 102.105 97.810 104.090 ;
        RECT 98.450 102.105 98.640 104.090 ;
        RECT 101.620 107.365 101.810 109.350 ;
        RECT 101.620 102.870 101.810 104.855 ;
        RECT 107.970 108.250 108.140 110.130 ;
        RECT 111.140 108.250 111.310 110.130 ;
        RECT 111.730 108.250 111.900 110.130 ;
        RECT 113.020 108.250 113.190 110.130 ;
        RECT 113.610 108.250 113.780 110.130 ;
        RECT 114.900 108.250 115.070 110.130 ;
        RECT 116.780 108.250 116.950 110.130 ;
        RECT 118.660 108.250 118.830 110.130 ;
        RECT 120.540 108.250 120.710 110.130 ;
        RECT 108.280 107.830 109.120 108.000 ;
        RECT 110.160 107.830 111.000 108.000 ;
        RECT 112.040 107.830 112.880 108.000 ;
        RECT 113.920 107.830 114.760 108.000 ;
        RECT 115.800 107.830 116.640 108.000 ;
        RECT 117.680 107.830 118.520 108.000 ;
        RECT 119.560 107.830 120.400 108.000 ;
        RECT 108.280 107.290 109.120 107.460 ;
        RECT 110.160 107.290 111.000 107.460 ;
        RECT 112.040 107.290 112.880 107.460 ;
        RECT 113.920 107.290 114.760 107.460 ;
        RECT 115.800 107.290 116.640 107.460 ;
        RECT 117.680 107.290 118.520 107.460 ;
        RECT 119.560 107.290 120.400 107.460 ;
        RECT 107.970 105.160 108.140 107.040 ;
        RECT 104.310 104.990 104.650 105.160 ;
        RECT 105.710 104.990 106.050 105.160 ;
        RECT 111.140 105.160 111.310 107.040 ;
        RECT 111.730 105.160 111.900 107.040 ;
        RECT 113.020 105.160 113.190 107.040 ;
        RECT 113.610 105.160 113.780 107.040 ;
        RECT 114.900 105.160 115.070 107.040 ;
        RECT 116.780 105.160 116.950 107.040 ;
        RECT 118.660 105.160 118.830 107.040 ;
        RECT 120.540 105.160 120.710 107.040 ;
        RECT 104.000 104.360 104.170 104.740 ;
        RECT 108.280 104.740 109.120 104.910 ;
        RECT 110.160 104.740 111.000 104.910 ;
        RECT 112.040 104.740 112.880 104.910 ;
        RECT 113.920 104.740 114.760 104.910 ;
        RECT 115.800 104.740 116.640 104.910 ;
        RECT 117.680 104.740 118.520 104.910 ;
        RECT 119.560 104.740 120.400 104.910 ;
        RECT 105.400 104.360 105.570 104.740 ;
        RECT 108.280 104.185 109.120 104.355 ;
        RECT 110.160 104.185 111.000 104.355 ;
        RECT 112.040 104.185 112.880 104.355 ;
        RECT 113.920 104.185 114.760 104.355 ;
        RECT 115.800 104.185 116.640 104.355 ;
        RECT 117.680 104.185 118.520 104.355 ;
        RECT 104.310 103.940 104.650 104.110 ;
        RECT 105.710 103.940 106.050 104.110 ;
        RECT 104.310 103.375 104.650 103.545 ;
        RECT 105.710 103.375 106.050 103.545 ;
        RECT 85.620 99.545 86.460 99.715 ;
        RECT 87.500 99.545 88.340 99.715 ;
        RECT 89.380 99.545 90.220 99.715 ;
        RECT 91.260 99.545 92.100 99.715 ;
        RECT 93.140 99.545 93.980 99.715 ;
        RECT 95.020 99.545 95.860 99.715 ;
        RECT 85.620 99.005 86.460 99.175 ;
        RECT 87.500 99.005 88.340 99.175 ;
        RECT 89.380 99.005 90.220 99.175 ;
        RECT 91.260 99.005 92.100 99.175 ;
        RECT 93.140 99.005 93.980 99.175 ;
        RECT 95.020 99.005 95.860 99.175 ;
        RECT 85.310 94.830 85.480 98.710 ;
        RECT 86.600 94.830 86.770 98.710 ;
        RECT 87.190 94.830 87.360 98.710 ;
        RECT 88.480 94.830 88.650 98.710 ;
        RECT 89.070 94.830 89.240 98.710 ;
        RECT 92.240 94.830 92.410 98.710 ;
        RECT 94.120 94.830 94.290 98.710 ;
        RECT 96.000 94.830 96.170 98.710 ;
        RECT 85.620 94.365 86.460 94.535 ;
        RECT 87.500 94.365 88.340 94.535 ;
        RECT 89.380 94.365 90.220 94.535 ;
        RECT 91.260 94.365 92.100 94.535 ;
        RECT 93.140 94.365 93.980 94.535 ;
        RECT 95.020 94.365 95.860 94.535 ;
        RECT 96.790 93.860 96.980 95.845 ;
        RECT 97.620 93.860 97.810 95.845 ;
        RECT 98.450 93.860 98.640 95.845 ;
        RECT 99.280 93.860 99.470 95.845 ;
        RECT 101.620 99.575 101.810 101.560 ;
        RECT 101.620 95.080 101.810 97.065 ;
        RECT 104.000 102.200 104.170 103.080 ;
        RECT 105.400 102.200 105.570 103.080 ;
        RECT 104.310 101.735 104.650 101.905 ;
        RECT 105.710 101.735 106.050 101.905 ;
        RECT 107.970 100.010 108.140 103.890 ;
        RECT 109.260 100.010 109.430 103.890 ;
        RECT 109.850 100.010 110.020 103.890 ;
        RECT 111.140 100.010 111.310 103.890 ;
        RECT 111.730 100.010 111.900 103.890 ;
        RECT 114.900 100.010 115.070 103.890 ;
        RECT 116.780 100.010 116.950 103.890 ;
        RECT 118.660 100.010 118.830 103.890 ;
        RECT 119.450 102.105 119.640 104.090 ;
        RECT 120.280 102.105 120.470 104.090 ;
        RECT 121.110 102.105 121.300 104.090 ;
        RECT 124.280 107.365 124.470 109.350 ;
        RECT 124.280 102.870 124.470 104.855 ;
        RECT 108.280 99.545 109.120 99.715 ;
        RECT 110.160 99.545 111.000 99.715 ;
        RECT 112.040 99.545 112.880 99.715 ;
        RECT 113.920 99.545 114.760 99.715 ;
        RECT 115.800 99.545 116.640 99.715 ;
        RECT 117.680 99.545 118.520 99.715 ;
        RECT 108.280 99.005 109.120 99.175 ;
        RECT 110.160 99.005 111.000 99.175 ;
        RECT 112.040 99.005 112.880 99.175 ;
        RECT 113.920 99.005 114.760 99.175 ;
        RECT 115.800 99.005 116.640 99.175 ;
        RECT 117.680 99.005 118.520 99.175 ;
        RECT 107.970 94.830 108.140 98.710 ;
        RECT 109.260 94.830 109.430 98.710 ;
        RECT 109.850 94.830 110.020 98.710 ;
        RECT 111.140 94.830 111.310 98.710 ;
        RECT 111.730 94.830 111.900 98.710 ;
        RECT 114.900 94.830 115.070 98.710 ;
        RECT 116.780 94.830 116.950 98.710 ;
        RECT 118.660 94.830 118.830 98.710 ;
        RECT 108.280 94.365 109.120 94.535 ;
        RECT 110.160 94.365 111.000 94.535 ;
        RECT 112.040 94.365 112.880 94.535 ;
        RECT 113.920 94.365 114.760 94.535 ;
        RECT 115.800 94.365 116.640 94.535 ;
        RECT 117.680 94.365 118.520 94.535 ;
        RECT 119.450 93.860 119.640 95.845 ;
        RECT 120.280 93.860 120.470 95.845 ;
        RECT 121.110 93.860 121.300 95.845 ;
        RECT 121.940 93.860 122.130 95.845 ;
        RECT 124.280 99.575 124.470 101.560 ;
        RECT 124.280 95.080 124.470 97.065 ;
        RECT 40.300 93.040 41.140 93.210 ;
        RECT 42.180 93.040 43.020 93.210 ;
        RECT 44.060 93.040 44.900 93.210 ;
        RECT 45.940 93.040 46.780 93.210 ;
        RECT 47.820 93.040 48.660 93.210 ;
        RECT 49.700 93.040 50.540 93.210 ;
        RECT 51.580 93.040 52.420 93.210 ;
        RECT 62.960 93.040 63.800 93.210 ;
        RECT 64.840 93.040 65.680 93.210 ;
        RECT 66.720 93.040 67.560 93.210 ;
        RECT 68.600 93.040 69.440 93.210 ;
        RECT 70.480 93.040 71.320 93.210 ;
        RECT 72.360 93.040 73.200 93.210 ;
        RECT 74.240 93.040 75.080 93.210 ;
        RECT 85.620 93.040 86.460 93.210 ;
        RECT 87.500 93.040 88.340 93.210 ;
        RECT 89.380 93.040 90.220 93.210 ;
        RECT 91.260 93.040 92.100 93.210 ;
        RECT 93.140 93.040 93.980 93.210 ;
        RECT 95.020 93.040 95.860 93.210 ;
        RECT 96.900 93.040 97.740 93.210 ;
        RECT 108.280 93.040 109.120 93.210 ;
        RECT 110.160 93.040 111.000 93.210 ;
        RECT 112.040 93.040 112.880 93.210 ;
        RECT 113.920 93.040 114.760 93.210 ;
        RECT 115.800 93.040 116.640 93.210 ;
        RECT 117.680 93.040 118.520 93.210 ;
        RECT 119.560 93.040 120.400 93.210 ;
        RECT 39.990 90.910 40.160 92.790 ;
        RECT 43.160 90.910 43.330 92.790 ;
        RECT 43.750 90.910 43.920 92.790 ;
        RECT 45.040 90.910 45.210 92.790 ;
        RECT 45.630 90.910 45.800 92.790 ;
        RECT 46.920 90.910 47.090 92.790 ;
        RECT 48.800 90.910 48.970 92.790 ;
        RECT 50.680 90.910 50.850 92.790 ;
        RECT 52.560 90.910 52.730 92.790 ;
        RECT 40.300 90.490 41.140 90.660 ;
        RECT 42.180 90.490 43.020 90.660 ;
        RECT 44.060 90.490 44.900 90.660 ;
        RECT 45.940 90.490 46.780 90.660 ;
        RECT 47.820 90.490 48.660 90.660 ;
        RECT 49.700 90.490 50.540 90.660 ;
        RECT 51.580 90.490 52.420 90.660 ;
        RECT 40.300 89.950 41.140 90.120 ;
        RECT 42.180 89.950 43.020 90.120 ;
        RECT 44.060 89.950 44.900 90.120 ;
        RECT 45.940 89.950 46.780 90.120 ;
        RECT 47.820 89.950 48.660 90.120 ;
        RECT 49.700 89.950 50.540 90.120 ;
        RECT 51.580 89.950 52.420 90.120 ;
        RECT 39.990 87.820 40.160 89.700 ;
        RECT 36.330 87.650 36.670 87.820 ;
        RECT 37.730 87.650 38.070 87.820 ;
        RECT 43.160 87.820 43.330 89.700 ;
        RECT 43.750 87.820 43.920 89.700 ;
        RECT 45.040 87.820 45.210 89.700 ;
        RECT 45.630 87.820 45.800 89.700 ;
        RECT 46.920 87.820 47.090 89.700 ;
        RECT 48.800 87.820 48.970 89.700 ;
        RECT 50.680 87.820 50.850 89.700 ;
        RECT 52.560 87.820 52.730 89.700 ;
        RECT 36.020 87.020 36.190 87.400 ;
        RECT 40.300 87.400 41.140 87.570 ;
        RECT 42.180 87.400 43.020 87.570 ;
        RECT 44.060 87.400 44.900 87.570 ;
        RECT 45.940 87.400 46.780 87.570 ;
        RECT 47.820 87.400 48.660 87.570 ;
        RECT 49.700 87.400 50.540 87.570 ;
        RECT 51.580 87.400 52.420 87.570 ;
        RECT 37.420 87.020 37.590 87.400 ;
        RECT 40.300 86.845 41.140 87.015 ;
        RECT 42.180 86.845 43.020 87.015 ;
        RECT 44.060 86.845 44.900 87.015 ;
        RECT 45.940 86.845 46.780 87.015 ;
        RECT 47.820 86.845 48.660 87.015 ;
        RECT 49.700 86.845 50.540 87.015 ;
        RECT 36.330 86.600 36.670 86.770 ;
        RECT 37.730 86.600 38.070 86.770 ;
        RECT 36.330 86.035 36.670 86.205 ;
        RECT 37.730 86.035 38.070 86.205 ;
        RECT 36.020 84.860 36.190 85.740 ;
        RECT 37.420 84.860 37.590 85.740 ;
        RECT 36.330 84.395 36.670 84.565 ;
        RECT 37.730 84.395 38.070 84.565 ;
        RECT 39.990 82.670 40.160 86.550 ;
        RECT 41.280 82.670 41.450 86.550 ;
        RECT 41.870 82.670 42.040 86.550 ;
        RECT 43.160 82.670 43.330 86.550 ;
        RECT 43.750 82.670 43.920 86.550 ;
        RECT 46.920 82.670 47.090 86.550 ;
        RECT 48.800 82.670 48.970 86.550 ;
        RECT 50.680 82.670 50.850 86.550 ;
        RECT 51.470 84.765 51.660 86.750 ;
        RECT 52.300 84.765 52.490 86.750 ;
        RECT 53.130 84.765 53.320 86.750 ;
        RECT 56.300 90.025 56.490 92.010 ;
        RECT 56.300 85.530 56.490 87.515 ;
        RECT 62.650 90.910 62.820 92.790 ;
        RECT 65.820 90.910 65.990 92.790 ;
        RECT 66.410 90.910 66.580 92.790 ;
        RECT 67.700 90.910 67.870 92.790 ;
        RECT 68.290 90.910 68.460 92.790 ;
        RECT 69.580 90.910 69.750 92.790 ;
        RECT 71.460 90.910 71.630 92.790 ;
        RECT 73.340 90.910 73.510 92.790 ;
        RECT 75.220 90.910 75.390 92.790 ;
        RECT 62.960 90.490 63.800 90.660 ;
        RECT 64.840 90.490 65.680 90.660 ;
        RECT 66.720 90.490 67.560 90.660 ;
        RECT 68.600 90.490 69.440 90.660 ;
        RECT 70.480 90.490 71.320 90.660 ;
        RECT 72.360 90.490 73.200 90.660 ;
        RECT 74.240 90.490 75.080 90.660 ;
        RECT 62.960 89.950 63.800 90.120 ;
        RECT 64.840 89.950 65.680 90.120 ;
        RECT 66.720 89.950 67.560 90.120 ;
        RECT 68.600 89.950 69.440 90.120 ;
        RECT 70.480 89.950 71.320 90.120 ;
        RECT 72.360 89.950 73.200 90.120 ;
        RECT 74.240 89.950 75.080 90.120 ;
        RECT 62.650 87.820 62.820 89.700 ;
        RECT 58.990 87.650 59.330 87.820 ;
        RECT 60.390 87.650 60.730 87.820 ;
        RECT 65.820 87.820 65.990 89.700 ;
        RECT 66.410 87.820 66.580 89.700 ;
        RECT 67.700 87.820 67.870 89.700 ;
        RECT 68.290 87.820 68.460 89.700 ;
        RECT 69.580 87.820 69.750 89.700 ;
        RECT 71.460 87.820 71.630 89.700 ;
        RECT 73.340 87.820 73.510 89.700 ;
        RECT 75.220 87.820 75.390 89.700 ;
        RECT 58.680 87.020 58.850 87.400 ;
        RECT 62.960 87.400 63.800 87.570 ;
        RECT 64.840 87.400 65.680 87.570 ;
        RECT 66.720 87.400 67.560 87.570 ;
        RECT 68.600 87.400 69.440 87.570 ;
        RECT 70.480 87.400 71.320 87.570 ;
        RECT 72.360 87.400 73.200 87.570 ;
        RECT 74.240 87.400 75.080 87.570 ;
        RECT 60.080 87.020 60.250 87.400 ;
        RECT 62.960 86.845 63.800 87.015 ;
        RECT 64.840 86.845 65.680 87.015 ;
        RECT 66.720 86.845 67.560 87.015 ;
        RECT 68.600 86.845 69.440 87.015 ;
        RECT 70.480 86.845 71.320 87.015 ;
        RECT 72.360 86.845 73.200 87.015 ;
        RECT 58.990 86.600 59.330 86.770 ;
        RECT 60.390 86.600 60.730 86.770 ;
        RECT 58.990 86.035 59.330 86.205 ;
        RECT 60.390 86.035 60.730 86.205 ;
        RECT 40.300 82.205 41.140 82.375 ;
        RECT 42.180 82.205 43.020 82.375 ;
        RECT 44.060 82.205 44.900 82.375 ;
        RECT 45.940 82.205 46.780 82.375 ;
        RECT 47.820 82.205 48.660 82.375 ;
        RECT 49.700 82.205 50.540 82.375 ;
        RECT 40.300 81.665 41.140 81.835 ;
        RECT 42.180 81.665 43.020 81.835 ;
        RECT 44.060 81.665 44.900 81.835 ;
        RECT 45.940 81.665 46.780 81.835 ;
        RECT 47.820 81.665 48.660 81.835 ;
        RECT 49.700 81.665 50.540 81.835 ;
        RECT 39.990 77.490 40.160 81.370 ;
        RECT 41.280 77.490 41.450 81.370 ;
        RECT 41.870 77.490 42.040 81.370 ;
        RECT 43.160 77.490 43.330 81.370 ;
        RECT 43.750 77.490 43.920 81.370 ;
        RECT 46.920 77.490 47.090 81.370 ;
        RECT 48.800 77.490 48.970 81.370 ;
        RECT 50.680 77.490 50.850 81.370 ;
        RECT 40.300 77.025 41.140 77.195 ;
        RECT 42.180 77.025 43.020 77.195 ;
        RECT 44.060 77.025 44.900 77.195 ;
        RECT 45.940 77.025 46.780 77.195 ;
        RECT 47.820 77.025 48.660 77.195 ;
        RECT 49.700 77.025 50.540 77.195 ;
        RECT 51.470 76.520 51.660 78.505 ;
        RECT 52.300 76.520 52.490 78.505 ;
        RECT 53.130 76.520 53.320 78.505 ;
        RECT 53.960 76.520 54.150 78.505 ;
        RECT 56.300 82.235 56.490 84.220 ;
        RECT 56.300 77.740 56.490 79.725 ;
        RECT 58.680 84.860 58.850 85.740 ;
        RECT 60.080 84.860 60.250 85.740 ;
        RECT 58.990 84.395 59.330 84.565 ;
        RECT 60.390 84.395 60.730 84.565 ;
        RECT 62.650 82.670 62.820 86.550 ;
        RECT 63.940 82.670 64.110 86.550 ;
        RECT 64.530 82.670 64.700 86.550 ;
        RECT 65.820 82.670 65.990 86.550 ;
        RECT 66.410 82.670 66.580 86.550 ;
        RECT 69.580 82.670 69.750 86.550 ;
        RECT 71.460 82.670 71.630 86.550 ;
        RECT 73.340 82.670 73.510 86.550 ;
        RECT 74.130 84.765 74.320 86.750 ;
        RECT 74.960 84.765 75.150 86.750 ;
        RECT 75.790 84.765 75.980 86.750 ;
        RECT 78.960 90.025 79.150 92.010 ;
        RECT 78.960 85.530 79.150 87.515 ;
        RECT 85.310 90.910 85.480 92.790 ;
        RECT 88.480 90.910 88.650 92.790 ;
        RECT 89.070 90.910 89.240 92.790 ;
        RECT 90.360 90.910 90.530 92.790 ;
        RECT 90.950 90.910 91.120 92.790 ;
        RECT 92.240 90.910 92.410 92.790 ;
        RECT 94.120 90.910 94.290 92.790 ;
        RECT 96.000 90.910 96.170 92.790 ;
        RECT 97.880 90.910 98.050 92.790 ;
        RECT 85.620 90.490 86.460 90.660 ;
        RECT 87.500 90.490 88.340 90.660 ;
        RECT 89.380 90.490 90.220 90.660 ;
        RECT 91.260 90.490 92.100 90.660 ;
        RECT 93.140 90.490 93.980 90.660 ;
        RECT 95.020 90.490 95.860 90.660 ;
        RECT 96.900 90.490 97.740 90.660 ;
        RECT 85.620 89.950 86.460 90.120 ;
        RECT 87.500 89.950 88.340 90.120 ;
        RECT 89.380 89.950 90.220 90.120 ;
        RECT 91.260 89.950 92.100 90.120 ;
        RECT 93.140 89.950 93.980 90.120 ;
        RECT 95.020 89.950 95.860 90.120 ;
        RECT 96.900 89.950 97.740 90.120 ;
        RECT 85.310 87.820 85.480 89.700 ;
        RECT 81.650 87.650 81.990 87.820 ;
        RECT 83.050 87.650 83.390 87.820 ;
        RECT 88.480 87.820 88.650 89.700 ;
        RECT 89.070 87.820 89.240 89.700 ;
        RECT 90.360 87.820 90.530 89.700 ;
        RECT 90.950 87.820 91.120 89.700 ;
        RECT 92.240 87.820 92.410 89.700 ;
        RECT 94.120 87.820 94.290 89.700 ;
        RECT 96.000 87.820 96.170 89.700 ;
        RECT 97.880 87.820 98.050 89.700 ;
        RECT 81.340 87.020 81.510 87.400 ;
        RECT 85.620 87.400 86.460 87.570 ;
        RECT 87.500 87.400 88.340 87.570 ;
        RECT 89.380 87.400 90.220 87.570 ;
        RECT 91.260 87.400 92.100 87.570 ;
        RECT 93.140 87.400 93.980 87.570 ;
        RECT 95.020 87.400 95.860 87.570 ;
        RECT 96.900 87.400 97.740 87.570 ;
        RECT 82.740 87.020 82.910 87.400 ;
        RECT 85.620 86.845 86.460 87.015 ;
        RECT 87.500 86.845 88.340 87.015 ;
        RECT 89.380 86.845 90.220 87.015 ;
        RECT 91.260 86.845 92.100 87.015 ;
        RECT 93.140 86.845 93.980 87.015 ;
        RECT 95.020 86.845 95.860 87.015 ;
        RECT 81.650 86.600 81.990 86.770 ;
        RECT 83.050 86.600 83.390 86.770 ;
        RECT 81.650 86.035 81.990 86.205 ;
        RECT 83.050 86.035 83.390 86.205 ;
        RECT 62.960 82.205 63.800 82.375 ;
        RECT 64.840 82.205 65.680 82.375 ;
        RECT 66.720 82.205 67.560 82.375 ;
        RECT 68.600 82.205 69.440 82.375 ;
        RECT 70.480 82.205 71.320 82.375 ;
        RECT 72.360 82.205 73.200 82.375 ;
        RECT 62.960 81.665 63.800 81.835 ;
        RECT 64.840 81.665 65.680 81.835 ;
        RECT 66.720 81.665 67.560 81.835 ;
        RECT 68.600 81.665 69.440 81.835 ;
        RECT 70.480 81.665 71.320 81.835 ;
        RECT 72.360 81.665 73.200 81.835 ;
        RECT 62.650 77.490 62.820 81.370 ;
        RECT 63.940 77.490 64.110 81.370 ;
        RECT 64.530 77.490 64.700 81.370 ;
        RECT 65.820 77.490 65.990 81.370 ;
        RECT 66.410 77.490 66.580 81.370 ;
        RECT 69.580 77.490 69.750 81.370 ;
        RECT 71.460 77.490 71.630 81.370 ;
        RECT 73.340 77.490 73.510 81.370 ;
        RECT 62.960 77.025 63.800 77.195 ;
        RECT 64.840 77.025 65.680 77.195 ;
        RECT 66.720 77.025 67.560 77.195 ;
        RECT 68.600 77.025 69.440 77.195 ;
        RECT 70.480 77.025 71.320 77.195 ;
        RECT 72.360 77.025 73.200 77.195 ;
        RECT 74.130 76.520 74.320 78.505 ;
        RECT 74.960 76.520 75.150 78.505 ;
        RECT 75.790 76.520 75.980 78.505 ;
        RECT 76.620 76.520 76.810 78.505 ;
        RECT 78.960 82.235 79.150 84.220 ;
        RECT 78.960 77.740 79.150 79.725 ;
        RECT 81.340 84.860 81.510 85.740 ;
        RECT 82.740 84.860 82.910 85.740 ;
        RECT 81.650 84.395 81.990 84.565 ;
        RECT 83.050 84.395 83.390 84.565 ;
        RECT 85.310 82.670 85.480 86.550 ;
        RECT 86.600 82.670 86.770 86.550 ;
        RECT 87.190 82.670 87.360 86.550 ;
        RECT 88.480 82.670 88.650 86.550 ;
        RECT 89.070 82.670 89.240 86.550 ;
        RECT 92.240 82.670 92.410 86.550 ;
        RECT 94.120 82.670 94.290 86.550 ;
        RECT 96.000 82.670 96.170 86.550 ;
        RECT 96.790 84.765 96.980 86.750 ;
        RECT 97.620 84.765 97.810 86.750 ;
        RECT 98.450 84.765 98.640 86.750 ;
        RECT 101.620 90.025 101.810 92.010 ;
        RECT 101.620 85.530 101.810 87.515 ;
        RECT 107.970 90.910 108.140 92.790 ;
        RECT 111.140 90.910 111.310 92.790 ;
        RECT 111.730 90.910 111.900 92.790 ;
        RECT 113.020 90.910 113.190 92.790 ;
        RECT 113.610 90.910 113.780 92.790 ;
        RECT 114.900 90.910 115.070 92.790 ;
        RECT 116.780 90.910 116.950 92.790 ;
        RECT 118.660 90.910 118.830 92.790 ;
        RECT 120.540 90.910 120.710 92.790 ;
        RECT 108.280 90.490 109.120 90.660 ;
        RECT 110.160 90.490 111.000 90.660 ;
        RECT 112.040 90.490 112.880 90.660 ;
        RECT 113.920 90.490 114.760 90.660 ;
        RECT 115.800 90.490 116.640 90.660 ;
        RECT 117.680 90.490 118.520 90.660 ;
        RECT 119.560 90.490 120.400 90.660 ;
        RECT 108.280 89.950 109.120 90.120 ;
        RECT 110.160 89.950 111.000 90.120 ;
        RECT 112.040 89.950 112.880 90.120 ;
        RECT 113.920 89.950 114.760 90.120 ;
        RECT 115.800 89.950 116.640 90.120 ;
        RECT 117.680 89.950 118.520 90.120 ;
        RECT 119.560 89.950 120.400 90.120 ;
        RECT 107.970 87.820 108.140 89.700 ;
        RECT 104.310 87.650 104.650 87.820 ;
        RECT 105.710 87.650 106.050 87.820 ;
        RECT 111.140 87.820 111.310 89.700 ;
        RECT 111.730 87.820 111.900 89.700 ;
        RECT 113.020 87.820 113.190 89.700 ;
        RECT 113.610 87.820 113.780 89.700 ;
        RECT 114.900 87.820 115.070 89.700 ;
        RECT 116.780 87.820 116.950 89.700 ;
        RECT 118.660 87.820 118.830 89.700 ;
        RECT 120.540 87.820 120.710 89.700 ;
        RECT 104.000 87.020 104.170 87.400 ;
        RECT 108.280 87.400 109.120 87.570 ;
        RECT 110.160 87.400 111.000 87.570 ;
        RECT 112.040 87.400 112.880 87.570 ;
        RECT 113.920 87.400 114.760 87.570 ;
        RECT 115.800 87.400 116.640 87.570 ;
        RECT 117.680 87.400 118.520 87.570 ;
        RECT 119.560 87.400 120.400 87.570 ;
        RECT 105.400 87.020 105.570 87.400 ;
        RECT 108.280 86.845 109.120 87.015 ;
        RECT 110.160 86.845 111.000 87.015 ;
        RECT 112.040 86.845 112.880 87.015 ;
        RECT 113.920 86.845 114.760 87.015 ;
        RECT 115.800 86.845 116.640 87.015 ;
        RECT 117.680 86.845 118.520 87.015 ;
        RECT 104.310 86.600 104.650 86.770 ;
        RECT 105.710 86.600 106.050 86.770 ;
        RECT 104.310 86.035 104.650 86.205 ;
        RECT 105.710 86.035 106.050 86.205 ;
        RECT 85.620 82.205 86.460 82.375 ;
        RECT 87.500 82.205 88.340 82.375 ;
        RECT 89.380 82.205 90.220 82.375 ;
        RECT 91.260 82.205 92.100 82.375 ;
        RECT 93.140 82.205 93.980 82.375 ;
        RECT 95.020 82.205 95.860 82.375 ;
        RECT 85.620 81.665 86.460 81.835 ;
        RECT 87.500 81.665 88.340 81.835 ;
        RECT 89.380 81.665 90.220 81.835 ;
        RECT 91.260 81.665 92.100 81.835 ;
        RECT 93.140 81.665 93.980 81.835 ;
        RECT 95.020 81.665 95.860 81.835 ;
        RECT 85.310 77.490 85.480 81.370 ;
        RECT 86.600 77.490 86.770 81.370 ;
        RECT 87.190 77.490 87.360 81.370 ;
        RECT 88.480 77.490 88.650 81.370 ;
        RECT 89.070 77.490 89.240 81.370 ;
        RECT 92.240 77.490 92.410 81.370 ;
        RECT 94.120 77.490 94.290 81.370 ;
        RECT 96.000 77.490 96.170 81.370 ;
        RECT 85.620 77.025 86.460 77.195 ;
        RECT 87.500 77.025 88.340 77.195 ;
        RECT 89.380 77.025 90.220 77.195 ;
        RECT 91.260 77.025 92.100 77.195 ;
        RECT 93.140 77.025 93.980 77.195 ;
        RECT 95.020 77.025 95.860 77.195 ;
        RECT 96.790 76.520 96.980 78.505 ;
        RECT 97.620 76.520 97.810 78.505 ;
        RECT 98.450 76.520 98.640 78.505 ;
        RECT 99.280 76.520 99.470 78.505 ;
        RECT 101.620 82.235 101.810 84.220 ;
        RECT 101.620 77.740 101.810 79.725 ;
        RECT 104.000 84.860 104.170 85.740 ;
        RECT 105.400 84.860 105.570 85.740 ;
        RECT 104.310 84.395 104.650 84.565 ;
        RECT 105.710 84.395 106.050 84.565 ;
        RECT 107.970 82.670 108.140 86.550 ;
        RECT 109.260 82.670 109.430 86.550 ;
        RECT 109.850 82.670 110.020 86.550 ;
        RECT 111.140 82.670 111.310 86.550 ;
        RECT 111.730 82.670 111.900 86.550 ;
        RECT 114.900 82.670 115.070 86.550 ;
        RECT 116.780 82.670 116.950 86.550 ;
        RECT 118.660 82.670 118.830 86.550 ;
        RECT 119.450 84.765 119.640 86.750 ;
        RECT 120.280 84.765 120.470 86.750 ;
        RECT 121.110 84.765 121.300 86.750 ;
        RECT 124.280 90.025 124.470 92.010 ;
        RECT 124.280 85.530 124.470 87.515 ;
        RECT 108.280 82.205 109.120 82.375 ;
        RECT 110.160 82.205 111.000 82.375 ;
        RECT 112.040 82.205 112.880 82.375 ;
        RECT 113.920 82.205 114.760 82.375 ;
        RECT 115.800 82.205 116.640 82.375 ;
        RECT 117.680 82.205 118.520 82.375 ;
        RECT 108.280 81.665 109.120 81.835 ;
        RECT 110.160 81.665 111.000 81.835 ;
        RECT 112.040 81.665 112.880 81.835 ;
        RECT 113.920 81.665 114.760 81.835 ;
        RECT 115.800 81.665 116.640 81.835 ;
        RECT 117.680 81.665 118.520 81.835 ;
        RECT 107.970 77.490 108.140 81.370 ;
        RECT 109.260 77.490 109.430 81.370 ;
        RECT 109.850 77.490 110.020 81.370 ;
        RECT 111.140 77.490 111.310 81.370 ;
        RECT 111.730 77.490 111.900 81.370 ;
        RECT 114.900 77.490 115.070 81.370 ;
        RECT 116.780 77.490 116.950 81.370 ;
        RECT 118.660 77.490 118.830 81.370 ;
        RECT 108.280 77.025 109.120 77.195 ;
        RECT 110.160 77.025 111.000 77.195 ;
        RECT 112.040 77.025 112.880 77.195 ;
        RECT 113.920 77.025 114.760 77.195 ;
        RECT 115.800 77.025 116.640 77.195 ;
        RECT 117.680 77.025 118.520 77.195 ;
        RECT 119.450 76.520 119.640 78.505 ;
        RECT 120.280 76.520 120.470 78.505 ;
        RECT 121.110 76.520 121.300 78.505 ;
        RECT 121.940 76.520 122.130 78.505 ;
        RECT 124.280 82.235 124.470 84.220 ;
        RECT 124.280 77.740 124.470 79.725 ;
        RECT 40.300 75.700 41.140 75.870 ;
        RECT 42.180 75.700 43.020 75.870 ;
        RECT 44.060 75.700 44.900 75.870 ;
        RECT 45.940 75.700 46.780 75.870 ;
        RECT 47.820 75.700 48.660 75.870 ;
        RECT 49.700 75.700 50.540 75.870 ;
        RECT 51.580 75.700 52.420 75.870 ;
        RECT 62.960 75.700 63.800 75.870 ;
        RECT 64.840 75.700 65.680 75.870 ;
        RECT 66.720 75.700 67.560 75.870 ;
        RECT 68.600 75.700 69.440 75.870 ;
        RECT 70.480 75.700 71.320 75.870 ;
        RECT 72.360 75.700 73.200 75.870 ;
        RECT 74.240 75.700 75.080 75.870 ;
        RECT 85.620 75.700 86.460 75.870 ;
        RECT 87.500 75.700 88.340 75.870 ;
        RECT 89.380 75.700 90.220 75.870 ;
        RECT 91.260 75.700 92.100 75.870 ;
        RECT 93.140 75.700 93.980 75.870 ;
        RECT 95.020 75.700 95.860 75.870 ;
        RECT 96.900 75.700 97.740 75.870 ;
        RECT 108.280 75.700 109.120 75.870 ;
        RECT 110.160 75.700 111.000 75.870 ;
        RECT 112.040 75.700 112.880 75.870 ;
        RECT 113.920 75.700 114.760 75.870 ;
        RECT 115.800 75.700 116.640 75.870 ;
        RECT 117.680 75.700 118.520 75.870 ;
        RECT 119.560 75.700 120.400 75.870 ;
        RECT 39.990 73.570 40.160 75.450 ;
        RECT 43.160 73.570 43.330 75.450 ;
        RECT 43.750 73.570 43.920 75.450 ;
        RECT 45.040 73.570 45.210 75.450 ;
        RECT 45.630 73.570 45.800 75.450 ;
        RECT 46.920 73.570 47.090 75.450 ;
        RECT 48.800 73.570 48.970 75.450 ;
        RECT 50.680 73.570 50.850 75.450 ;
        RECT 52.560 73.570 52.730 75.450 ;
        RECT 40.300 73.150 41.140 73.320 ;
        RECT 42.180 73.150 43.020 73.320 ;
        RECT 44.060 73.150 44.900 73.320 ;
        RECT 45.940 73.150 46.780 73.320 ;
        RECT 47.820 73.150 48.660 73.320 ;
        RECT 49.700 73.150 50.540 73.320 ;
        RECT 51.580 73.150 52.420 73.320 ;
        RECT 40.300 72.610 41.140 72.780 ;
        RECT 42.180 72.610 43.020 72.780 ;
        RECT 44.060 72.610 44.900 72.780 ;
        RECT 45.940 72.610 46.780 72.780 ;
        RECT 47.820 72.610 48.660 72.780 ;
        RECT 49.700 72.610 50.540 72.780 ;
        RECT 51.580 72.610 52.420 72.780 ;
        RECT 39.990 70.480 40.160 72.360 ;
        RECT 36.330 70.310 36.670 70.480 ;
        RECT 37.730 70.310 38.070 70.480 ;
        RECT 43.160 70.480 43.330 72.360 ;
        RECT 43.750 70.480 43.920 72.360 ;
        RECT 45.040 70.480 45.210 72.360 ;
        RECT 45.630 70.480 45.800 72.360 ;
        RECT 46.920 70.480 47.090 72.360 ;
        RECT 48.800 70.480 48.970 72.360 ;
        RECT 50.680 70.480 50.850 72.360 ;
        RECT 52.560 70.480 52.730 72.360 ;
        RECT 36.020 69.680 36.190 70.060 ;
        RECT 40.300 70.060 41.140 70.230 ;
        RECT 42.180 70.060 43.020 70.230 ;
        RECT 44.060 70.060 44.900 70.230 ;
        RECT 45.940 70.060 46.780 70.230 ;
        RECT 47.820 70.060 48.660 70.230 ;
        RECT 49.700 70.060 50.540 70.230 ;
        RECT 51.580 70.060 52.420 70.230 ;
        RECT 37.420 69.680 37.590 70.060 ;
        RECT 40.300 69.505 41.140 69.675 ;
        RECT 42.180 69.505 43.020 69.675 ;
        RECT 44.060 69.505 44.900 69.675 ;
        RECT 45.940 69.505 46.780 69.675 ;
        RECT 47.820 69.505 48.660 69.675 ;
        RECT 49.700 69.505 50.540 69.675 ;
        RECT 36.330 69.260 36.670 69.430 ;
        RECT 37.730 69.260 38.070 69.430 ;
        RECT 36.330 68.695 36.670 68.865 ;
        RECT 37.730 68.695 38.070 68.865 ;
        RECT 36.020 67.520 36.190 68.400 ;
        RECT 37.420 67.520 37.590 68.400 ;
        RECT 36.330 67.055 36.670 67.225 ;
        RECT 37.730 67.055 38.070 67.225 ;
        RECT 39.990 65.330 40.160 69.210 ;
        RECT 41.280 65.330 41.450 69.210 ;
        RECT 41.870 65.330 42.040 69.210 ;
        RECT 43.160 65.330 43.330 69.210 ;
        RECT 43.750 65.330 43.920 69.210 ;
        RECT 46.920 65.330 47.090 69.210 ;
        RECT 48.800 65.330 48.970 69.210 ;
        RECT 50.680 65.330 50.850 69.210 ;
        RECT 51.470 67.425 51.660 69.410 ;
        RECT 52.300 67.425 52.490 69.410 ;
        RECT 53.130 67.425 53.320 69.410 ;
        RECT 56.300 72.685 56.490 74.670 ;
        RECT 56.300 68.190 56.490 70.175 ;
        RECT 62.650 73.570 62.820 75.450 ;
        RECT 65.820 73.570 65.990 75.450 ;
        RECT 66.410 73.570 66.580 75.450 ;
        RECT 67.700 73.570 67.870 75.450 ;
        RECT 68.290 73.570 68.460 75.450 ;
        RECT 69.580 73.570 69.750 75.450 ;
        RECT 71.460 73.570 71.630 75.450 ;
        RECT 73.340 73.570 73.510 75.450 ;
        RECT 75.220 73.570 75.390 75.450 ;
        RECT 62.960 73.150 63.800 73.320 ;
        RECT 64.840 73.150 65.680 73.320 ;
        RECT 66.720 73.150 67.560 73.320 ;
        RECT 68.600 73.150 69.440 73.320 ;
        RECT 70.480 73.150 71.320 73.320 ;
        RECT 72.360 73.150 73.200 73.320 ;
        RECT 74.240 73.150 75.080 73.320 ;
        RECT 62.960 72.610 63.800 72.780 ;
        RECT 64.840 72.610 65.680 72.780 ;
        RECT 66.720 72.610 67.560 72.780 ;
        RECT 68.600 72.610 69.440 72.780 ;
        RECT 70.480 72.610 71.320 72.780 ;
        RECT 72.360 72.610 73.200 72.780 ;
        RECT 74.240 72.610 75.080 72.780 ;
        RECT 62.650 70.480 62.820 72.360 ;
        RECT 58.990 70.310 59.330 70.480 ;
        RECT 60.390 70.310 60.730 70.480 ;
        RECT 65.820 70.480 65.990 72.360 ;
        RECT 66.410 70.480 66.580 72.360 ;
        RECT 67.700 70.480 67.870 72.360 ;
        RECT 68.290 70.480 68.460 72.360 ;
        RECT 69.580 70.480 69.750 72.360 ;
        RECT 71.460 70.480 71.630 72.360 ;
        RECT 73.340 70.480 73.510 72.360 ;
        RECT 75.220 70.480 75.390 72.360 ;
        RECT 58.680 69.680 58.850 70.060 ;
        RECT 62.960 70.060 63.800 70.230 ;
        RECT 64.840 70.060 65.680 70.230 ;
        RECT 66.720 70.060 67.560 70.230 ;
        RECT 68.600 70.060 69.440 70.230 ;
        RECT 70.480 70.060 71.320 70.230 ;
        RECT 72.360 70.060 73.200 70.230 ;
        RECT 74.240 70.060 75.080 70.230 ;
        RECT 60.080 69.680 60.250 70.060 ;
        RECT 62.960 69.505 63.800 69.675 ;
        RECT 64.840 69.505 65.680 69.675 ;
        RECT 66.720 69.505 67.560 69.675 ;
        RECT 68.600 69.505 69.440 69.675 ;
        RECT 70.480 69.505 71.320 69.675 ;
        RECT 72.360 69.505 73.200 69.675 ;
        RECT 58.990 69.260 59.330 69.430 ;
        RECT 60.390 69.260 60.730 69.430 ;
        RECT 58.990 68.695 59.330 68.865 ;
        RECT 60.390 68.695 60.730 68.865 ;
        RECT 40.300 64.865 41.140 65.035 ;
        RECT 42.180 64.865 43.020 65.035 ;
        RECT 44.060 64.865 44.900 65.035 ;
        RECT 45.940 64.865 46.780 65.035 ;
        RECT 47.820 64.865 48.660 65.035 ;
        RECT 49.700 64.865 50.540 65.035 ;
        RECT 40.300 64.325 41.140 64.495 ;
        RECT 42.180 64.325 43.020 64.495 ;
        RECT 44.060 64.325 44.900 64.495 ;
        RECT 45.940 64.325 46.780 64.495 ;
        RECT 47.820 64.325 48.660 64.495 ;
        RECT 49.700 64.325 50.540 64.495 ;
        RECT 39.990 60.150 40.160 64.030 ;
        RECT 41.280 60.150 41.450 64.030 ;
        RECT 41.870 60.150 42.040 64.030 ;
        RECT 43.160 60.150 43.330 64.030 ;
        RECT 43.750 60.150 43.920 64.030 ;
        RECT 46.920 60.150 47.090 64.030 ;
        RECT 48.800 60.150 48.970 64.030 ;
        RECT 50.680 60.150 50.850 64.030 ;
        RECT 40.300 59.685 41.140 59.855 ;
        RECT 42.180 59.685 43.020 59.855 ;
        RECT 44.060 59.685 44.900 59.855 ;
        RECT 45.940 59.685 46.780 59.855 ;
        RECT 47.820 59.685 48.660 59.855 ;
        RECT 49.700 59.685 50.540 59.855 ;
        RECT 51.470 59.180 51.660 61.165 ;
        RECT 52.300 59.180 52.490 61.165 ;
        RECT 53.130 59.180 53.320 61.165 ;
        RECT 53.960 59.180 54.150 61.165 ;
        RECT 56.300 64.895 56.490 66.880 ;
        RECT 56.300 60.400 56.490 62.385 ;
        RECT 58.680 67.520 58.850 68.400 ;
        RECT 60.080 67.520 60.250 68.400 ;
        RECT 58.990 67.055 59.330 67.225 ;
        RECT 60.390 67.055 60.730 67.225 ;
        RECT 62.650 65.330 62.820 69.210 ;
        RECT 63.940 65.330 64.110 69.210 ;
        RECT 64.530 65.330 64.700 69.210 ;
        RECT 65.820 65.330 65.990 69.210 ;
        RECT 66.410 65.330 66.580 69.210 ;
        RECT 69.580 65.330 69.750 69.210 ;
        RECT 71.460 65.330 71.630 69.210 ;
        RECT 73.340 65.330 73.510 69.210 ;
        RECT 74.130 67.425 74.320 69.410 ;
        RECT 74.960 67.425 75.150 69.410 ;
        RECT 75.790 67.425 75.980 69.410 ;
        RECT 78.960 72.685 79.150 74.670 ;
        RECT 78.960 68.190 79.150 70.175 ;
        RECT 85.310 73.570 85.480 75.450 ;
        RECT 88.480 73.570 88.650 75.450 ;
        RECT 89.070 73.570 89.240 75.450 ;
        RECT 90.360 73.570 90.530 75.450 ;
        RECT 90.950 73.570 91.120 75.450 ;
        RECT 92.240 73.570 92.410 75.450 ;
        RECT 94.120 73.570 94.290 75.450 ;
        RECT 96.000 73.570 96.170 75.450 ;
        RECT 97.880 73.570 98.050 75.450 ;
        RECT 85.620 73.150 86.460 73.320 ;
        RECT 87.500 73.150 88.340 73.320 ;
        RECT 89.380 73.150 90.220 73.320 ;
        RECT 91.260 73.150 92.100 73.320 ;
        RECT 93.140 73.150 93.980 73.320 ;
        RECT 95.020 73.150 95.860 73.320 ;
        RECT 96.900 73.150 97.740 73.320 ;
        RECT 85.620 72.610 86.460 72.780 ;
        RECT 87.500 72.610 88.340 72.780 ;
        RECT 89.380 72.610 90.220 72.780 ;
        RECT 91.260 72.610 92.100 72.780 ;
        RECT 93.140 72.610 93.980 72.780 ;
        RECT 95.020 72.610 95.860 72.780 ;
        RECT 96.900 72.610 97.740 72.780 ;
        RECT 85.310 70.480 85.480 72.360 ;
        RECT 81.650 70.310 81.990 70.480 ;
        RECT 83.050 70.310 83.390 70.480 ;
        RECT 88.480 70.480 88.650 72.360 ;
        RECT 89.070 70.480 89.240 72.360 ;
        RECT 90.360 70.480 90.530 72.360 ;
        RECT 90.950 70.480 91.120 72.360 ;
        RECT 92.240 70.480 92.410 72.360 ;
        RECT 94.120 70.480 94.290 72.360 ;
        RECT 96.000 70.480 96.170 72.360 ;
        RECT 97.880 70.480 98.050 72.360 ;
        RECT 81.340 69.680 81.510 70.060 ;
        RECT 85.620 70.060 86.460 70.230 ;
        RECT 87.500 70.060 88.340 70.230 ;
        RECT 89.380 70.060 90.220 70.230 ;
        RECT 91.260 70.060 92.100 70.230 ;
        RECT 93.140 70.060 93.980 70.230 ;
        RECT 95.020 70.060 95.860 70.230 ;
        RECT 96.900 70.060 97.740 70.230 ;
        RECT 82.740 69.680 82.910 70.060 ;
        RECT 85.620 69.505 86.460 69.675 ;
        RECT 87.500 69.505 88.340 69.675 ;
        RECT 89.380 69.505 90.220 69.675 ;
        RECT 91.260 69.505 92.100 69.675 ;
        RECT 93.140 69.505 93.980 69.675 ;
        RECT 95.020 69.505 95.860 69.675 ;
        RECT 81.650 69.260 81.990 69.430 ;
        RECT 83.050 69.260 83.390 69.430 ;
        RECT 81.650 68.695 81.990 68.865 ;
        RECT 83.050 68.695 83.390 68.865 ;
        RECT 62.960 64.865 63.800 65.035 ;
        RECT 64.840 64.865 65.680 65.035 ;
        RECT 66.720 64.865 67.560 65.035 ;
        RECT 68.600 64.865 69.440 65.035 ;
        RECT 70.480 64.865 71.320 65.035 ;
        RECT 72.360 64.865 73.200 65.035 ;
        RECT 62.960 64.325 63.800 64.495 ;
        RECT 64.840 64.325 65.680 64.495 ;
        RECT 66.720 64.325 67.560 64.495 ;
        RECT 68.600 64.325 69.440 64.495 ;
        RECT 70.480 64.325 71.320 64.495 ;
        RECT 72.360 64.325 73.200 64.495 ;
        RECT 62.650 60.150 62.820 64.030 ;
        RECT 63.940 60.150 64.110 64.030 ;
        RECT 64.530 60.150 64.700 64.030 ;
        RECT 65.820 60.150 65.990 64.030 ;
        RECT 66.410 60.150 66.580 64.030 ;
        RECT 69.580 60.150 69.750 64.030 ;
        RECT 71.460 60.150 71.630 64.030 ;
        RECT 73.340 60.150 73.510 64.030 ;
        RECT 62.960 59.685 63.800 59.855 ;
        RECT 64.840 59.685 65.680 59.855 ;
        RECT 66.720 59.685 67.560 59.855 ;
        RECT 68.600 59.685 69.440 59.855 ;
        RECT 70.480 59.685 71.320 59.855 ;
        RECT 72.360 59.685 73.200 59.855 ;
        RECT 74.130 59.180 74.320 61.165 ;
        RECT 74.960 59.180 75.150 61.165 ;
        RECT 75.790 59.180 75.980 61.165 ;
        RECT 76.620 59.180 76.810 61.165 ;
        RECT 78.960 64.895 79.150 66.880 ;
        RECT 78.960 60.400 79.150 62.385 ;
        RECT 81.340 67.520 81.510 68.400 ;
        RECT 82.740 67.520 82.910 68.400 ;
        RECT 81.650 67.055 81.990 67.225 ;
        RECT 83.050 67.055 83.390 67.225 ;
        RECT 85.310 65.330 85.480 69.210 ;
        RECT 86.600 65.330 86.770 69.210 ;
        RECT 87.190 65.330 87.360 69.210 ;
        RECT 88.480 65.330 88.650 69.210 ;
        RECT 89.070 65.330 89.240 69.210 ;
        RECT 92.240 65.330 92.410 69.210 ;
        RECT 94.120 65.330 94.290 69.210 ;
        RECT 96.000 65.330 96.170 69.210 ;
        RECT 96.790 67.425 96.980 69.410 ;
        RECT 97.620 67.425 97.810 69.410 ;
        RECT 98.450 67.425 98.640 69.410 ;
        RECT 101.620 72.685 101.810 74.670 ;
        RECT 101.620 68.190 101.810 70.175 ;
        RECT 107.970 73.570 108.140 75.450 ;
        RECT 111.140 73.570 111.310 75.450 ;
        RECT 111.730 73.570 111.900 75.450 ;
        RECT 113.020 73.570 113.190 75.450 ;
        RECT 113.610 73.570 113.780 75.450 ;
        RECT 114.900 73.570 115.070 75.450 ;
        RECT 116.780 73.570 116.950 75.450 ;
        RECT 118.660 73.570 118.830 75.450 ;
        RECT 120.540 73.570 120.710 75.450 ;
        RECT 108.280 73.150 109.120 73.320 ;
        RECT 110.160 73.150 111.000 73.320 ;
        RECT 112.040 73.150 112.880 73.320 ;
        RECT 113.920 73.150 114.760 73.320 ;
        RECT 115.800 73.150 116.640 73.320 ;
        RECT 117.680 73.150 118.520 73.320 ;
        RECT 119.560 73.150 120.400 73.320 ;
        RECT 108.280 72.610 109.120 72.780 ;
        RECT 110.160 72.610 111.000 72.780 ;
        RECT 112.040 72.610 112.880 72.780 ;
        RECT 113.920 72.610 114.760 72.780 ;
        RECT 115.800 72.610 116.640 72.780 ;
        RECT 117.680 72.610 118.520 72.780 ;
        RECT 119.560 72.610 120.400 72.780 ;
        RECT 107.970 70.480 108.140 72.360 ;
        RECT 104.310 70.310 104.650 70.480 ;
        RECT 105.710 70.310 106.050 70.480 ;
        RECT 111.140 70.480 111.310 72.360 ;
        RECT 111.730 70.480 111.900 72.360 ;
        RECT 113.020 70.480 113.190 72.360 ;
        RECT 113.610 70.480 113.780 72.360 ;
        RECT 114.900 70.480 115.070 72.360 ;
        RECT 116.780 70.480 116.950 72.360 ;
        RECT 118.660 70.480 118.830 72.360 ;
        RECT 120.540 70.480 120.710 72.360 ;
        RECT 104.000 69.680 104.170 70.060 ;
        RECT 108.280 70.060 109.120 70.230 ;
        RECT 110.160 70.060 111.000 70.230 ;
        RECT 112.040 70.060 112.880 70.230 ;
        RECT 113.920 70.060 114.760 70.230 ;
        RECT 115.800 70.060 116.640 70.230 ;
        RECT 117.680 70.060 118.520 70.230 ;
        RECT 119.560 70.060 120.400 70.230 ;
        RECT 105.400 69.680 105.570 70.060 ;
        RECT 108.280 69.505 109.120 69.675 ;
        RECT 110.160 69.505 111.000 69.675 ;
        RECT 112.040 69.505 112.880 69.675 ;
        RECT 113.920 69.505 114.760 69.675 ;
        RECT 115.800 69.505 116.640 69.675 ;
        RECT 117.680 69.505 118.520 69.675 ;
        RECT 104.310 69.260 104.650 69.430 ;
        RECT 105.710 69.260 106.050 69.430 ;
        RECT 104.310 68.695 104.650 68.865 ;
        RECT 105.710 68.695 106.050 68.865 ;
        RECT 85.620 64.865 86.460 65.035 ;
        RECT 87.500 64.865 88.340 65.035 ;
        RECT 89.380 64.865 90.220 65.035 ;
        RECT 91.260 64.865 92.100 65.035 ;
        RECT 93.140 64.865 93.980 65.035 ;
        RECT 95.020 64.865 95.860 65.035 ;
        RECT 85.620 64.325 86.460 64.495 ;
        RECT 87.500 64.325 88.340 64.495 ;
        RECT 89.380 64.325 90.220 64.495 ;
        RECT 91.260 64.325 92.100 64.495 ;
        RECT 93.140 64.325 93.980 64.495 ;
        RECT 95.020 64.325 95.860 64.495 ;
        RECT 85.310 60.150 85.480 64.030 ;
        RECT 86.600 60.150 86.770 64.030 ;
        RECT 87.190 60.150 87.360 64.030 ;
        RECT 88.480 60.150 88.650 64.030 ;
        RECT 89.070 60.150 89.240 64.030 ;
        RECT 92.240 60.150 92.410 64.030 ;
        RECT 94.120 60.150 94.290 64.030 ;
        RECT 96.000 60.150 96.170 64.030 ;
        RECT 85.620 59.685 86.460 59.855 ;
        RECT 87.500 59.685 88.340 59.855 ;
        RECT 89.380 59.685 90.220 59.855 ;
        RECT 91.260 59.685 92.100 59.855 ;
        RECT 93.140 59.685 93.980 59.855 ;
        RECT 95.020 59.685 95.860 59.855 ;
        RECT 96.790 59.180 96.980 61.165 ;
        RECT 97.620 59.180 97.810 61.165 ;
        RECT 98.450 59.180 98.640 61.165 ;
        RECT 99.280 59.180 99.470 61.165 ;
        RECT 101.620 64.895 101.810 66.880 ;
        RECT 101.620 60.400 101.810 62.385 ;
        RECT 104.000 67.520 104.170 68.400 ;
        RECT 105.400 67.520 105.570 68.400 ;
        RECT 104.310 67.055 104.650 67.225 ;
        RECT 105.710 67.055 106.050 67.225 ;
        RECT 107.970 65.330 108.140 69.210 ;
        RECT 109.260 65.330 109.430 69.210 ;
        RECT 109.850 65.330 110.020 69.210 ;
        RECT 111.140 65.330 111.310 69.210 ;
        RECT 111.730 65.330 111.900 69.210 ;
        RECT 114.900 65.330 115.070 69.210 ;
        RECT 116.780 65.330 116.950 69.210 ;
        RECT 118.660 65.330 118.830 69.210 ;
        RECT 119.450 67.425 119.640 69.410 ;
        RECT 120.280 67.425 120.470 69.410 ;
        RECT 121.110 67.425 121.300 69.410 ;
        RECT 124.280 72.685 124.470 74.670 ;
        RECT 124.280 68.190 124.470 70.175 ;
        RECT 108.280 64.865 109.120 65.035 ;
        RECT 110.160 64.865 111.000 65.035 ;
        RECT 112.040 64.865 112.880 65.035 ;
        RECT 113.920 64.865 114.760 65.035 ;
        RECT 115.800 64.865 116.640 65.035 ;
        RECT 117.680 64.865 118.520 65.035 ;
        RECT 108.280 64.325 109.120 64.495 ;
        RECT 110.160 64.325 111.000 64.495 ;
        RECT 112.040 64.325 112.880 64.495 ;
        RECT 113.920 64.325 114.760 64.495 ;
        RECT 115.800 64.325 116.640 64.495 ;
        RECT 117.680 64.325 118.520 64.495 ;
        RECT 107.970 60.150 108.140 64.030 ;
        RECT 109.260 60.150 109.430 64.030 ;
        RECT 109.850 60.150 110.020 64.030 ;
        RECT 111.140 60.150 111.310 64.030 ;
        RECT 111.730 60.150 111.900 64.030 ;
        RECT 114.900 60.150 115.070 64.030 ;
        RECT 116.780 60.150 116.950 64.030 ;
        RECT 118.660 60.150 118.830 64.030 ;
        RECT 108.280 59.685 109.120 59.855 ;
        RECT 110.160 59.685 111.000 59.855 ;
        RECT 112.040 59.685 112.880 59.855 ;
        RECT 113.920 59.685 114.760 59.855 ;
        RECT 115.800 59.685 116.640 59.855 ;
        RECT 117.680 59.685 118.520 59.855 ;
        RECT 119.450 59.180 119.640 61.165 ;
        RECT 120.280 59.180 120.470 61.165 ;
        RECT 121.110 59.180 121.300 61.165 ;
        RECT 121.940 59.180 122.130 61.165 ;
        RECT 124.280 64.895 124.470 66.880 ;
        RECT 124.280 60.400 124.470 62.385 ;
        RECT 40.300 57.700 41.140 57.870 ;
        RECT 42.180 57.700 43.020 57.870 ;
        RECT 44.060 57.700 44.900 57.870 ;
        RECT 47.820 57.700 48.660 57.870 ;
        RECT 49.700 57.700 50.540 57.870 ;
        RECT 51.580 57.700 52.420 57.870 ;
        RECT 62.960 57.700 63.800 57.870 ;
        RECT 64.840 57.700 65.680 57.870 ;
        RECT 66.720 57.700 67.560 57.870 ;
        RECT 70.480 57.700 71.320 57.870 ;
        RECT 72.360 57.700 73.200 57.870 ;
        RECT 74.240 57.700 75.080 57.870 ;
        RECT 85.620 57.700 86.460 57.870 ;
        RECT 87.500 57.700 88.340 57.870 ;
        RECT 89.380 57.700 90.220 57.870 ;
        RECT 93.140 57.700 93.980 57.870 ;
        RECT 95.020 57.700 95.860 57.870 ;
        RECT 96.900 57.700 97.740 57.870 ;
        RECT 108.280 57.700 109.120 57.870 ;
        RECT 110.160 57.700 111.000 57.870 ;
        RECT 112.040 57.700 112.880 57.870 ;
        RECT 115.800 57.700 116.640 57.870 ;
        RECT 117.680 57.700 118.520 57.870 ;
        RECT 119.560 57.700 120.400 57.870 ;
        RECT 39.990 55.570 40.160 57.450 ;
        RECT 43.160 55.570 43.330 57.450 ;
        RECT 43.750 55.570 43.920 57.450 ;
        RECT 45.040 55.570 45.210 57.450 ;
        RECT 45.630 55.570 45.800 57.450 ;
        RECT 46.920 55.570 47.090 57.450 ;
        RECT 48.800 55.570 48.970 57.450 ;
        RECT 50.680 55.570 50.850 57.450 ;
        RECT 52.560 55.570 52.730 57.450 ;
        RECT 62.650 55.570 62.820 57.450 ;
        RECT 65.820 55.570 65.990 57.450 ;
        RECT 66.410 55.570 66.580 57.450 ;
        RECT 67.700 55.570 67.870 57.450 ;
        RECT 68.290 55.570 68.460 57.450 ;
        RECT 69.580 55.570 69.750 57.450 ;
        RECT 71.460 55.570 71.630 57.450 ;
        RECT 73.340 55.570 73.510 57.450 ;
        RECT 75.220 55.570 75.390 57.450 ;
        RECT 85.310 55.570 85.480 57.450 ;
        RECT 88.480 55.570 88.650 57.450 ;
        RECT 89.070 55.570 89.240 57.450 ;
        RECT 90.360 55.570 90.530 57.450 ;
        RECT 90.950 55.570 91.120 57.450 ;
        RECT 92.240 55.570 92.410 57.450 ;
        RECT 94.120 55.570 94.290 57.450 ;
        RECT 96.000 55.570 96.170 57.450 ;
        RECT 97.880 55.570 98.050 57.450 ;
        RECT 107.970 55.570 108.140 57.450 ;
        RECT 111.140 55.570 111.310 57.450 ;
        RECT 111.730 55.570 111.900 57.450 ;
        RECT 113.020 55.570 113.190 57.450 ;
        RECT 113.610 55.570 113.780 57.450 ;
        RECT 114.900 55.570 115.070 57.450 ;
        RECT 116.780 55.570 116.950 57.450 ;
        RECT 118.660 55.570 118.830 57.450 ;
        RECT 120.540 55.570 120.710 57.450 ;
        RECT 40.300 55.150 41.140 55.320 ;
        RECT 42.180 55.150 43.020 55.320 ;
        RECT 44.060 55.150 44.900 55.320 ;
        RECT 47.820 55.150 48.660 55.320 ;
        RECT 49.700 55.150 50.540 55.320 ;
        RECT 51.580 55.150 52.420 55.320 ;
        RECT 62.960 55.150 63.800 55.320 ;
        RECT 64.840 55.150 65.680 55.320 ;
        RECT 66.720 55.150 67.560 55.320 ;
        RECT 70.480 55.150 71.320 55.320 ;
        RECT 72.360 55.150 73.200 55.320 ;
        RECT 74.240 55.150 75.080 55.320 ;
        RECT 85.620 55.150 86.460 55.320 ;
        RECT 87.500 55.150 88.340 55.320 ;
        RECT 89.380 55.150 90.220 55.320 ;
        RECT 93.140 55.150 93.980 55.320 ;
        RECT 95.020 55.150 95.860 55.320 ;
        RECT 96.900 55.150 97.740 55.320 ;
        RECT 108.280 55.150 109.120 55.320 ;
        RECT 110.160 55.150 111.000 55.320 ;
        RECT 112.040 55.150 112.880 55.320 ;
        RECT 115.800 55.150 116.640 55.320 ;
        RECT 117.680 55.150 118.520 55.320 ;
        RECT 119.560 55.150 120.400 55.320 ;
        RECT 40.300 54.610 41.140 54.780 ;
        RECT 42.180 54.610 43.020 54.780 ;
        RECT 44.060 54.610 44.900 54.780 ;
        RECT 47.820 54.610 48.660 54.780 ;
        RECT 49.700 54.610 50.540 54.780 ;
        RECT 51.580 54.610 52.420 54.780 ;
        RECT 62.960 54.610 63.800 54.780 ;
        RECT 64.840 54.610 65.680 54.780 ;
        RECT 66.720 54.610 67.560 54.780 ;
        RECT 70.480 54.610 71.320 54.780 ;
        RECT 72.360 54.610 73.200 54.780 ;
        RECT 74.240 54.610 75.080 54.780 ;
        RECT 85.620 54.610 86.460 54.780 ;
        RECT 87.500 54.610 88.340 54.780 ;
        RECT 89.380 54.610 90.220 54.780 ;
        RECT 93.140 54.610 93.980 54.780 ;
        RECT 95.020 54.610 95.860 54.780 ;
        RECT 96.900 54.610 97.740 54.780 ;
        RECT 108.280 54.610 109.120 54.780 ;
        RECT 110.160 54.610 111.000 54.780 ;
        RECT 112.040 54.610 112.880 54.780 ;
        RECT 115.800 54.610 116.640 54.780 ;
        RECT 117.680 54.610 118.520 54.780 ;
        RECT 119.560 54.610 120.400 54.780 ;
        RECT 39.990 52.480 40.160 54.360 ;
        RECT 43.160 52.480 43.330 54.360 ;
        RECT 43.750 52.480 43.920 54.360 ;
        RECT 45.040 52.480 45.210 54.360 ;
        RECT 45.630 52.480 45.800 54.360 ;
        RECT 46.920 52.480 47.090 54.360 ;
        RECT 48.800 52.480 48.970 54.360 ;
        RECT 50.680 52.480 50.850 54.360 ;
        RECT 52.560 52.480 52.730 54.360 ;
        RECT 62.650 52.480 62.820 54.360 ;
        RECT 65.820 52.480 65.990 54.360 ;
        RECT 66.410 52.480 66.580 54.360 ;
        RECT 67.700 52.480 67.870 54.360 ;
        RECT 68.290 52.480 68.460 54.360 ;
        RECT 69.580 52.480 69.750 54.360 ;
        RECT 71.460 52.480 71.630 54.360 ;
        RECT 73.340 52.480 73.510 54.360 ;
        RECT 75.220 52.480 75.390 54.360 ;
        RECT 85.310 52.480 85.480 54.360 ;
        RECT 88.480 52.480 88.650 54.360 ;
        RECT 89.070 52.480 89.240 54.360 ;
        RECT 90.360 52.480 90.530 54.360 ;
        RECT 90.950 52.480 91.120 54.360 ;
        RECT 92.240 52.480 92.410 54.360 ;
        RECT 94.120 52.480 94.290 54.360 ;
        RECT 96.000 52.480 96.170 54.360 ;
        RECT 97.880 52.480 98.050 54.360 ;
        RECT 107.970 52.480 108.140 54.360 ;
        RECT 111.140 52.480 111.310 54.360 ;
        RECT 111.730 52.480 111.900 54.360 ;
        RECT 113.020 52.480 113.190 54.360 ;
        RECT 113.610 52.480 113.780 54.360 ;
        RECT 114.900 52.480 115.070 54.360 ;
        RECT 116.780 52.480 116.950 54.360 ;
        RECT 118.660 52.480 118.830 54.360 ;
        RECT 120.540 52.480 120.710 54.360 ;
        RECT 40.300 52.060 41.140 52.230 ;
        RECT 42.180 52.060 43.020 52.230 ;
        RECT 44.060 52.060 44.900 52.230 ;
        RECT 47.820 52.060 48.660 52.230 ;
        RECT 49.700 52.060 50.540 52.230 ;
        RECT 51.580 52.060 52.420 52.230 ;
        RECT 62.960 52.060 63.800 52.230 ;
        RECT 64.840 52.060 65.680 52.230 ;
        RECT 66.720 52.060 67.560 52.230 ;
        RECT 70.480 52.060 71.320 52.230 ;
        RECT 72.360 52.060 73.200 52.230 ;
        RECT 74.240 52.060 75.080 52.230 ;
        RECT 85.620 52.060 86.460 52.230 ;
        RECT 87.500 52.060 88.340 52.230 ;
        RECT 89.380 52.060 90.220 52.230 ;
        RECT 93.140 52.060 93.980 52.230 ;
        RECT 95.020 52.060 95.860 52.230 ;
        RECT 96.900 52.060 97.740 52.230 ;
        RECT 108.280 52.060 109.120 52.230 ;
        RECT 110.160 52.060 111.000 52.230 ;
        RECT 112.040 52.060 112.880 52.230 ;
        RECT 115.800 52.060 116.640 52.230 ;
        RECT 117.680 52.060 118.520 52.230 ;
        RECT 119.560 52.060 120.400 52.230 ;
        RECT 40.300 51.505 41.140 51.675 ;
        RECT 44.060 51.505 44.900 51.675 ;
        RECT 45.940 51.505 46.780 51.675 ;
        RECT 47.820 51.505 48.660 51.675 ;
        RECT 49.700 51.505 50.540 51.675 ;
        RECT 62.960 51.505 63.800 51.675 ;
        RECT 66.720 51.505 67.560 51.675 ;
        RECT 68.600 51.505 69.440 51.675 ;
        RECT 70.480 51.505 71.320 51.675 ;
        RECT 72.360 51.505 73.200 51.675 ;
        RECT 85.620 51.505 86.460 51.675 ;
        RECT 89.380 51.505 90.220 51.675 ;
        RECT 91.260 51.505 92.100 51.675 ;
        RECT 93.140 51.505 93.980 51.675 ;
        RECT 95.020 51.505 95.860 51.675 ;
        RECT 108.280 51.505 109.120 51.675 ;
        RECT 112.040 51.505 112.880 51.675 ;
        RECT 113.920 51.505 114.760 51.675 ;
        RECT 115.800 51.505 116.640 51.675 ;
        RECT 117.680 51.505 118.520 51.675 ;
        RECT 39.990 47.330 40.160 51.210 ;
        RECT 41.280 47.330 41.450 51.210 ;
        RECT 41.870 47.330 42.040 51.210 ;
        RECT 43.160 47.330 43.330 51.210 ;
        RECT 43.750 47.330 43.920 51.210 ;
        RECT 46.920 47.330 47.090 51.210 ;
        RECT 48.800 47.330 48.970 51.210 ;
        RECT 50.680 47.330 50.850 51.210 ;
        RECT 51.470 49.425 51.660 51.410 ;
        RECT 52.300 49.425 52.490 51.410 ;
        RECT 53.130 49.425 53.320 51.410 ;
        RECT 62.650 47.330 62.820 51.210 ;
        RECT 63.940 47.330 64.110 51.210 ;
        RECT 64.530 47.330 64.700 51.210 ;
        RECT 65.820 47.330 65.990 51.210 ;
        RECT 66.410 47.330 66.580 51.210 ;
        RECT 69.580 47.330 69.750 51.210 ;
        RECT 71.460 47.330 71.630 51.210 ;
        RECT 73.340 47.330 73.510 51.210 ;
        RECT 74.130 49.425 74.320 51.410 ;
        RECT 74.960 49.425 75.150 51.410 ;
        RECT 75.790 49.425 75.980 51.410 ;
        RECT 85.310 47.330 85.480 51.210 ;
        RECT 86.600 47.330 86.770 51.210 ;
        RECT 87.190 47.330 87.360 51.210 ;
        RECT 88.480 47.330 88.650 51.210 ;
        RECT 89.070 47.330 89.240 51.210 ;
        RECT 92.240 47.330 92.410 51.210 ;
        RECT 94.120 47.330 94.290 51.210 ;
        RECT 96.000 47.330 96.170 51.210 ;
        RECT 96.790 49.425 96.980 51.410 ;
        RECT 97.620 49.425 97.810 51.410 ;
        RECT 98.450 49.425 98.640 51.410 ;
        RECT 107.970 47.330 108.140 51.210 ;
        RECT 109.260 47.330 109.430 51.210 ;
        RECT 109.850 47.330 110.020 51.210 ;
        RECT 111.140 47.330 111.310 51.210 ;
        RECT 111.730 47.330 111.900 51.210 ;
        RECT 114.900 47.330 115.070 51.210 ;
        RECT 116.780 47.330 116.950 51.210 ;
        RECT 118.660 47.330 118.830 51.210 ;
        RECT 119.450 49.425 119.640 51.410 ;
        RECT 120.280 49.425 120.470 51.410 ;
        RECT 121.110 49.425 121.300 51.410 ;
        RECT 40.300 46.865 41.140 47.035 ;
        RECT 44.060 46.865 44.900 47.035 ;
        RECT 45.940 46.865 46.780 47.035 ;
        RECT 47.820 46.865 48.660 47.035 ;
        RECT 49.700 46.865 50.540 47.035 ;
        RECT 62.960 46.865 63.800 47.035 ;
        RECT 66.720 46.865 67.560 47.035 ;
        RECT 68.600 46.865 69.440 47.035 ;
        RECT 70.480 46.865 71.320 47.035 ;
        RECT 72.360 46.865 73.200 47.035 ;
        RECT 85.620 46.865 86.460 47.035 ;
        RECT 89.380 46.865 90.220 47.035 ;
        RECT 91.260 46.865 92.100 47.035 ;
        RECT 93.140 46.865 93.980 47.035 ;
        RECT 95.020 46.865 95.860 47.035 ;
        RECT 108.280 46.865 109.120 47.035 ;
        RECT 112.040 46.865 112.880 47.035 ;
        RECT 113.920 46.865 114.760 47.035 ;
        RECT 115.800 46.865 116.640 47.035 ;
        RECT 117.680 46.865 118.520 47.035 ;
        RECT 40.300 46.325 41.140 46.495 ;
        RECT 44.060 46.325 44.900 46.495 ;
        RECT 45.940 46.325 46.780 46.495 ;
        RECT 47.820 46.325 48.660 46.495 ;
        RECT 49.700 46.325 50.540 46.495 ;
        RECT 62.960 46.325 63.800 46.495 ;
        RECT 66.720 46.325 67.560 46.495 ;
        RECT 68.600 46.325 69.440 46.495 ;
        RECT 70.480 46.325 71.320 46.495 ;
        RECT 72.360 46.325 73.200 46.495 ;
        RECT 85.620 46.325 86.460 46.495 ;
        RECT 89.380 46.325 90.220 46.495 ;
        RECT 91.260 46.325 92.100 46.495 ;
        RECT 93.140 46.325 93.980 46.495 ;
        RECT 95.020 46.325 95.860 46.495 ;
        RECT 108.280 46.325 109.120 46.495 ;
        RECT 112.040 46.325 112.880 46.495 ;
        RECT 113.920 46.325 114.760 46.495 ;
        RECT 115.800 46.325 116.640 46.495 ;
        RECT 117.680 46.325 118.520 46.495 ;
        RECT 39.990 42.150 40.160 46.030 ;
        RECT 41.280 42.150 41.450 46.030 ;
        RECT 41.870 42.150 42.040 46.030 ;
        RECT 43.160 42.150 43.330 46.030 ;
        RECT 43.750 42.150 43.920 46.030 ;
        RECT 46.920 42.150 47.090 46.030 ;
        RECT 48.800 42.150 48.970 46.030 ;
        RECT 50.680 42.150 50.850 46.030 ;
        RECT 40.300 41.685 41.140 41.855 ;
        RECT 44.060 41.685 44.900 41.855 ;
        RECT 45.940 41.685 46.780 41.855 ;
        RECT 47.820 41.685 48.660 41.855 ;
        RECT 49.700 41.685 50.540 41.855 ;
        RECT 51.470 41.180 51.660 43.165 ;
        RECT 52.300 41.180 52.490 43.165 ;
        RECT 53.130 41.180 53.320 43.165 ;
        RECT 53.960 41.180 54.150 43.165 ;
        RECT 62.650 42.150 62.820 46.030 ;
        RECT 63.940 42.150 64.110 46.030 ;
        RECT 64.530 42.150 64.700 46.030 ;
        RECT 65.820 42.150 65.990 46.030 ;
        RECT 66.410 42.150 66.580 46.030 ;
        RECT 69.580 42.150 69.750 46.030 ;
        RECT 71.460 42.150 71.630 46.030 ;
        RECT 73.340 42.150 73.510 46.030 ;
        RECT 62.960 41.685 63.800 41.855 ;
        RECT 66.720 41.685 67.560 41.855 ;
        RECT 68.600 41.685 69.440 41.855 ;
        RECT 70.480 41.685 71.320 41.855 ;
        RECT 72.360 41.685 73.200 41.855 ;
        RECT 74.130 41.180 74.320 43.165 ;
        RECT 74.960 41.180 75.150 43.165 ;
        RECT 75.790 41.180 75.980 43.165 ;
        RECT 76.620 41.180 76.810 43.165 ;
        RECT 85.310 42.150 85.480 46.030 ;
        RECT 86.600 42.150 86.770 46.030 ;
        RECT 87.190 42.150 87.360 46.030 ;
        RECT 88.480 42.150 88.650 46.030 ;
        RECT 89.070 42.150 89.240 46.030 ;
        RECT 92.240 42.150 92.410 46.030 ;
        RECT 94.120 42.150 94.290 46.030 ;
        RECT 96.000 42.150 96.170 46.030 ;
        RECT 85.620 41.685 86.460 41.855 ;
        RECT 89.380 41.685 90.220 41.855 ;
        RECT 91.260 41.685 92.100 41.855 ;
        RECT 93.140 41.685 93.980 41.855 ;
        RECT 95.020 41.685 95.860 41.855 ;
        RECT 96.790 41.180 96.980 43.165 ;
        RECT 97.620 41.180 97.810 43.165 ;
        RECT 98.450 41.180 98.640 43.165 ;
        RECT 99.280 41.180 99.470 43.165 ;
        RECT 107.970 42.150 108.140 46.030 ;
        RECT 109.260 42.150 109.430 46.030 ;
        RECT 109.850 42.150 110.020 46.030 ;
        RECT 111.140 42.150 111.310 46.030 ;
        RECT 111.730 42.150 111.900 46.030 ;
        RECT 114.900 42.150 115.070 46.030 ;
        RECT 116.780 42.150 116.950 46.030 ;
        RECT 118.660 42.150 118.830 46.030 ;
        RECT 108.280 41.685 109.120 41.855 ;
        RECT 112.040 41.685 112.880 41.855 ;
        RECT 113.920 41.685 114.760 41.855 ;
        RECT 115.800 41.685 116.640 41.855 ;
        RECT 117.680 41.685 118.520 41.855 ;
        RECT 119.450 41.180 119.640 43.165 ;
        RECT 120.280 41.180 120.470 43.165 ;
        RECT 121.110 41.180 121.300 43.165 ;
        RECT 121.940 41.180 122.130 43.165 ;
      LAYER met1 ;
        RECT 76.350 187.850 76.670 187.910 ;
        RECT 93.370 187.850 93.690 187.910 ;
        RECT 76.350 187.710 93.690 187.850 ;
        RECT 76.350 187.650 76.670 187.710 ;
        RECT 93.370 187.650 93.690 187.710 ;
        RECT 74.510 187.510 74.830 187.570 ;
        RECT 117.290 187.510 117.610 187.570 ;
        RECT 74.510 187.370 117.610 187.510 ;
        RECT 74.510 187.310 74.830 187.370 ;
        RECT 117.290 187.310 117.610 187.370 ;
        RECT 83.710 185.810 84.030 185.870 ;
        RECT 87.405 185.810 87.695 185.855 ;
        RECT 83.710 185.670 87.695 185.810 ;
        RECT 83.710 185.610 84.030 185.670 ;
        RECT 87.405 185.625 87.695 185.670 ;
        RECT 108.105 185.810 108.395 185.855 ;
        RECT 110.390 185.810 110.710 185.870 ;
        RECT 108.105 185.670 110.710 185.810 ;
        RECT 108.105 185.625 108.395 185.670 ;
        RECT 110.390 185.610 110.710 185.670 ;
        RECT 102.110 185.270 102.430 185.530 ;
        RECT 106.710 185.470 107.030 185.530 ;
        RECT 112.230 185.470 112.550 185.530 ;
        RECT 106.710 185.330 112.550 185.470 ;
        RECT 106.710 185.270 107.030 185.330 ;
        RECT 112.230 185.270 112.550 185.330 ;
        RECT 57.030 185.130 57.350 185.190 ;
        RECT 57.505 185.130 57.795 185.175 ;
        RECT 57.030 184.990 57.795 185.130 ;
        RECT 57.030 184.930 57.350 184.990 ;
        RECT 57.505 184.945 57.795 184.990 ;
        RECT 58.410 185.130 58.730 185.190 ;
        RECT 59.345 185.130 59.635 185.175 ;
        RECT 58.410 184.990 59.635 185.130 ;
        RECT 58.410 184.930 58.730 184.990 ;
        RECT 59.345 184.945 59.635 184.990 ;
        RECT 62.550 184.930 62.870 185.190 ;
        RECT 65.770 184.930 66.090 185.190 ;
        RECT 69.465 184.945 69.755 185.175 ;
        RECT 63.485 184.790 63.775 184.835 ;
        RECT 63.930 184.790 64.250 184.850 ;
        RECT 63.485 184.650 64.250 184.790 ;
        RECT 69.540 184.790 69.680 184.945 ;
        RECT 69.910 184.930 70.230 185.190 ;
        RECT 73.130 184.930 73.450 185.190 ;
        RECT 75.890 184.930 76.210 185.190 ;
        RECT 78.205 185.130 78.495 185.175 ;
        RECT 83.250 185.130 83.570 185.190 ;
        RECT 78.205 184.990 83.570 185.130 ;
        RECT 78.205 184.945 78.495 184.990 ;
        RECT 83.250 184.930 83.570 184.990 ;
        RECT 84.185 184.945 84.475 185.175 ;
        RECT 97.065 185.130 97.355 185.175 ;
        RECT 98.430 185.130 98.750 185.190 ;
        RECT 97.065 184.990 98.750 185.130 ;
        RECT 97.065 184.945 97.355 184.990 ;
        RECT 73.590 184.790 73.910 184.850 ;
        RECT 69.540 184.650 73.910 184.790 ;
        RECT 63.485 184.605 63.775 184.650 ;
        RECT 63.930 184.590 64.250 184.650 ;
        RECT 73.590 184.590 73.910 184.650 ;
        RECT 84.260 184.450 84.400 184.945 ;
        RECT 98.430 184.930 98.750 184.990 ;
        RECT 86.485 184.790 86.775 184.835 ;
        RECT 93.830 184.790 94.150 184.850 ;
        RECT 86.485 184.650 94.150 184.790 ;
        RECT 86.485 184.605 86.775 184.650 ;
        RECT 93.830 184.590 94.150 184.650 ;
        RECT 100.730 184.590 101.050 184.850 ;
        RECT 109.930 184.790 110.250 184.850 ;
        RECT 111.785 184.790 112.075 184.835 ;
        RECT 109.930 184.650 112.075 184.790 ;
        RECT 109.930 184.590 110.250 184.650 ;
        RECT 111.785 184.605 112.075 184.650 ;
        RECT 88.770 184.450 89.090 184.510 ;
        RECT 84.260 184.310 89.090 184.450 ;
        RECT 88.770 184.250 89.090 184.310 ;
        RECT 89.230 184.250 89.550 184.510 ;
        RECT 91.070 184.250 91.390 184.510 ;
        RECT 103.030 184.250 103.350 184.510 ;
        RECT 103.505 184.450 103.795 184.495 ;
        RECT 103.950 184.450 104.270 184.510 ;
        RECT 103.505 184.310 104.270 184.450 ;
        RECT 103.505 184.265 103.795 184.310 ;
        RECT 103.950 184.250 104.270 184.310 ;
        RECT 105.345 184.450 105.635 184.495 ;
        RECT 108.090 184.450 108.410 184.510 ;
        RECT 105.345 184.310 108.410 184.450 ;
        RECT 105.345 184.265 105.635 184.310 ;
        RECT 108.090 184.250 108.410 184.310 ;
        RECT 109.470 184.250 109.790 184.510 ;
        RECT 111.325 184.450 111.615 184.495 ;
        RECT 113.150 184.450 113.470 184.510 ;
        RECT 111.325 184.310 113.470 184.450 ;
        RECT 111.325 184.265 111.615 184.310 ;
        RECT 113.150 184.250 113.470 184.310 ;
        RECT 67.150 183.230 67.470 183.490 ;
        RECT 72.685 183.430 72.975 183.475 ;
        RECT 73.130 183.430 73.450 183.490 ;
        RECT 72.685 183.290 73.450 183.430 ;
        RECT 72.685 183.245 72.975 183.290 ;
        RECT 73.130 183.230 73.450 183.290 ;
        RECT 74.510 183.230 74.830 183.490 ;
        RECT 74.970 183.430 75.290 183.490 ;
        RECT 83.710 183.430 84.030 183.490 ;
        RECT 74.970 183.290 84.030 183.430 ;
        RECT 74.970 183.230 75.290 183.290 ;
        RECT 83.710 183.230 84.030 183.290 ;
        RECT 84.185 183.430 84.475 183.475 ;
        RECT 89.230 183.430 89.550 183.490 ;
        RECT 84.185 183.290 89.550 183.430 ;
        RECT 84.185 183.245 84.475 183.290 ;
        RECT 89.230 183.230 89.550 183.290 ;
        RECT 93.830 183.230 94.150 183.490 ;
        RECT 97.985 183.430 98.275 183.475 ;
        RECT 98.430 183.430 98.750 183.490 ;
        RECT 97.985 183.290 98.750 183.430 ;
        RECT 97.985 183.245 98.275 183.290 ;
        RECT 98.430 183.230 98.750 183.290 ;
        RECT 99.825 183.430 100.115 183.475 ;
        RECT 100.270 183.430 100.590 183.490 ;
        RECT 113.150 183.430 113.470 183.490 ;
        RECT 99.825 183.290 113.470 183.430 ;
        RECT 99.825 183.245 100.115 183.290 ;
        RECT 100.270 183.230 100.590 183.290 ;
        RECT 113.150 183.230 113.470 183.290 ;
        RECT 55.190 182.890 55.510 183.150 ;
        RECT 70.385 183.090 70.675 183.135 ;
        RECT 89.705 183.090 89.995 183.135 ;
        RECT 90.610 183.090 90.930 183.150 ;
        RECT 61.720 182.950 69.220 183.090 ;
        RECT 56.570 182.550 56.890 182.810 ;
        RECT 57.965 182.410 58.255 182.455 ;
        RECT 61.720 182.410 61.860 182.950 ;
        RECT 62.090 182.750 62.410 182.810 ;
        RECT 65.325 182.750 65.615 182.795 ;
        RECT 62.090 182.610 65.615 182.750 ;
        RECT 62.090 182.550 62.410 182.610 ;
        RECT 65.325 182.565 65.615 182.610 ;
        RECT 63.470 182.410 63.790 182.470 ;
        RECT 57.965 182.270 63.790 182.410 ;
        RECT 57.965 182.225 58.255 182.270 ;
        RECT 63.470 182.210 63.790 182.270 ;
        RECT 64.405 182.225 64.695 182.455 ;
        RECT 64.865 182.225 65.155 182.455 ;
        RECT 69.080 182.410 69.220 182.950 ;
        RECT 70.385 182.950 80.260 183.090 ;
        RECT 70.385 182.905 70.675 182.950 ;
        RECT 70.845 182.750 71.135 182.795 ;
        RECT 74.985 182.750 75.275 182.795 ;
        RECT 77.270 182.750 77.590 182.810 ;
        RECT 80.120 182.795 80.260 182.950 ;
        RECT 89.705 182.950 90.930 183.090 ;
        RECT 89.705 182.905 89.995 182.950 ;
        RECT 90.610 182.890 90.930 182.950 ;
        RECT 93.370 183.090 93.690 183.150 ;
        RECT 103.045 183.090 103.335 183.135 ;
        RECT 93.370 182.950 103.335 183.090 ;
        RECT 93.370 182.890 93.690 182.950 ;
        RECT 103.045 182.905 103.335 182.950 ;
        RECT 108.090 183.090 108.410 183.150 ;
        RECT 108.090 182.950 111.080 183.090 ;
        RECT 108.090 182.890 108.410 182.950 ;
        RECT 70.845 182.610 77.590 182.750 ;
        RECT 70.845 182.565 71.135 182.610 ;
        RECT 74.985 182.565 75.275 182.610 ;
        RECT 77.270 182.550 77.590 182.610 ;
        RECT 80.045 182.750 80.335 182.795 ;
        RECT 81.870 182.750 82.190 182.810 ;
        RECT 80.045 182.610 82.190 182.750 ;
        RECT 80.045 182.565 80.335 182.610 ;
        RECT 81.870 182.550 82.190 182.610 ;
        RECT 83.250 182.550 83.570 182.810 ;
        RECT 83.725 182.750 84.015 182.795 ;
        RECT 85.550 182.750 85.870 182.810 ;
        RECT 83.725 182.610 85.870 182.750 ;
        RECT 83.725 182.565 84.015 182.610 ;
        RECT 85.550 182.550 85.870 182.610 ;
        RECT 89.780 182.610 90.840 182.750 ;
        RECT 69.465 182.410 69.755 182.455 ;
        RECT 69.080 182.270 69.755 182.410 ;
        RECT 69.465 182.225 69.755 182.270 ;
        RECT 72.670 182.410 72.990 182.470 ;
        RECT 74.065 182.410 74.355 182.455 ;
        RECT 76.350 182.410 76.670 182.470 ;
        RECT 72.670 182.270 76.670 182.410 ;
        RECT 53.365 182.070 53.655 182.115 ;
        RECT 54.270 182.070 54.590 182.130 ;
        RECT 53.365 181.930 54.590 182.070 ;
        RECT 53.365 181.885 53.655 181.930 ;
        RECT 54.270 181.870 54.590 181.930 ;
        RECT 56.125 182.070 56.415 182.115 ;
        RECT 57.045 182.070 57.335 182.115 ;
        RECT 56.125 181.930 57.335 182.070 ;
        RECT 56.125 181.885 56.415 181.930 ;
        RECT 57.045 181.885 57.335 181.930 ;
        RECT 53.810 181.730 54.130 181.790 ;
        RECT 55.205 181.730 55.495 181.775 ;
        RECT 53.810 181.590 55.495 181.730 ;
        RECT 64.480 181.730 64.620 182.225 ;
        RECT 64.940 182.070 65.080 182.225 ;
        RECT 72.670 182.210 72.990 182.270 ;
        RECT 74.065 182.225 74.355 182.270 ;
        RECT 76.350 182.210 76.670 182.270 ;
        RECT 81.425 182.410 81.715 182.455 ;
        RECT 81.425 182.270 82.100 182.410 ;
        RECT 81.425 182.225 81.715 182.270 ;
        RECT 81.960 182.115 82.100 182.270 ;
        RECT 64.940 181.930 77.500 182.070 ;
        RECT 72.670 181.730 72.990 181.790 ;
        RECT 64.480 181.590 72.990 181.730 ;
        RECT 53.810 181.530 54.130 181.590 ;
        RECT 55.205 181.545 55.495 181.590 ;
        RECT 72.670 181.530 72.990 181.590 ;
        RECT 76.810 181.530 77.130 181.790 ;
        RECT 77.360 181.730 77.500 181.930 ;
        RECT 81.885 181.885 82.175 182.115 ;
        RECT 83.340 182.070 83.480 182.550 ;
        RECT 85.105 182.410 85.395 182.455 ;
        RECT 86.010 182.410 86.330 182.470 ;
        RECT 85.105 182.270 86.330 182.410 ;
        RECT 85.105 182.225 85.395 182.270 ;
        RECT 86.010 182.210 86.330 182.270 ;
        RECT 86.470 182.410 86.790 182.470 ;
        RECT 89.780 182.410 89.920 182.610 ;
        RECT 86.470 182.270 89.920 182.410 ;
        RECT 86.470 182.210 86.790 182.270 ;
        RECT 90.150 182.210 90.470 182.470 ;
        RECT 90.700 182.455 90.840 182.610 ;
        RECT 95.670 182.550 95.990 182.810 ;
        RECT 96.145 182.750 96.435 182.795 ;
        RECT 102.570 182.750 102.890 182.810 ;
        RECT 105.805 182.750 106.095 182.795 ;
        RECT 106.710 182.750 107.030 182.810 ;
        RECT 96.145 182.610 101.880 182.750 ;
        RECT 96.145 182.565 96.435 182.610 ;
        RECT 101.740 182.470 101.880 182.610 ;
        RECT 102.570 182.610 107.030 182.750 ;
        RECT 102.570 182.550 102.890 182.610 ;
        RECT 105.805 182.565 106.095 182.610 ;
        RECT 106.710 182.550 107.030 182.610 ;
        RECT 108.550 182.550 108.870 182.810 ;
        RECT 110.940 182.795 111.080 182.950 ;
        RECT 110.865 182.565 111.155 182.795 ;
        RECT 90.625 182.410 90.915 182.455 ;
        RECT 94.750 182.410 95.070 182.470 ;
        RECT 90.625 182.270 95.070 182.410 ;
        RECT 90.625 182.225 90.915 182.270 ;
        RECT 94.750 182.210 95.070 182.270 ;
        RECT 96.605 182.225 96.895 182.455 ;
        RECT 98.890 182.410 99.210 182.470 ;
        RECT 100.285 182.410 100.575 182.455 ;
        RECT 98.890 182.270 100.575 182.410 ;
        RECT 87.865 182.070 88.155 182.115 ;
        RECT 83.340 181.930 88.155 182.070 ;
        RECT 87.865 181.885 88.155 181.930 ;
        RECT 89.690 182.070 90.010 182.130 ;
        RECT 96.680 182.070 96.820 182.225 ;
        RECT 98.890 182.210 99.210 182.270 ;
        RECT 100.285 182.225 100.575 182.270 ;
        RECT 100.745 182.225 101.035 182.455 ;
        RECT 100.820 182.070 100.960 182.225 ;
        RECT 101.650 182.210 101.970 182.470 ;
        RECT 109.010 182.210 109.330 182.470 ;
        RECT 109.485 182.225 109.775 182.455 ;
        RECT 102.110 182.070 102.430 182.130 ;
        RECT 89.690 181.930 102.430 182.070 ;
        RECT 89.690 181.870 90.010 181.930 ;
        RECT 102.110 181.870 102.430 181.930 ;
        RECT 103.490 182.070 103.810 182.130 ;
        RECT 109.560 182.070 109.700 182.225 ;
        RECT 103.490 181.930 109.700 182.070 ;
        RECT 103.490 181.870 103.810 181.930 ;
        RECT 92.005 181.730 92.295 181.775 ;
        RECT 77.360 181.590 92.295 181.730 ;
        RECT 92.005 181.545 92.295 181.590 ;
        RECT 95.210 181.730 95.530 181.790 ;
        RECT 100.270 181.730 100.590 181.790 ;
        RECT 95.210 181.590 100.590 181.730 ;
        RECT 95.210 181.530 95.530 181.590 ;
        RECT 100.270 181.530 100.590 181.590 ;
        RECT 106.725 181.730 107.015 181.775 ;
        RECT 107.630 181.730 107.950 181.790 ;
        RECT 106.725 181.590 107.950 181.730 ;
        RECT 106.725 181.545 107.015 181.590 ;
        RECT 107.630 181.530 107.950 181.590 ;
        RECT 62.550 180.710 62.870 180.770 ;
        RECT 63.025 180.710 63.315 180.755 ;
        RECT 62.550 180.570 63.315 180.710 ;
        RECT 62.550 180.510 62.870 180.570 ;
        RECT 63.025 180.525 63.315 180.570 ;
        RECT 64.850 180.710 65.170 180.770 ;
        RECT 85.550 180.710 85.870 180.770 ;
        RECT 64.850 180.570 85.870 180.710 ;
        RECT 64.850 180.510 65.170 180.570 ;
        RECT 85.550 180.510 85.870 180.570 ;
        RECT 91.990 180.710 92.310 180.770 ;
        RECT 93.845 180.710 94.135 180.755 ;
        RECT 91.990 180.570 94.135 180.710 ;
        RECT 91.990 180.510 92.310 180.570 ;
        RECT 93.845 180.525 94.135 180.570 ;
        RECT 94.750 180.710 95.070 180.770 ;
        RECT 95.685 180.710 95.975 180.755 ;
        RECT 94.750 180.570 95.975 180.710 ;
        RECT 94.750 180.510 95.070 180.570 ;
        RECT 95.685 180.525 95.975 180.570 ;
        RECT 100.285 180.710 100.575 180.755 ;
        RECT 100.730 180.710 101.050 180.770 ;
        RECT 100.285 180.570 101.050 180.710 ;
        RECT 100.285 180.525 100.575 180.570 ;
        RECT 100.730 180.510 101.050 180.570 ;
        RECT 101.650 180.710 101.970 180.770 ;
        RECT 101.650 180.570 110.620 180.710 ;
        RECT 101.650 180.510 101.970 180.570 ;
        RECT 83.250 180.370 83.570 180.430 ;
        RECT 97.065 180.370 97.355 180.415 ;
        RECT 83.250 180.230 97.355 180.370 ;
        RECT 83.250 180.170 83.570 180.230 ;
        RECT 97.065 180.185 97.355 180.230 ;
        RECT 66.230 179.830 66.550 180.090 ;
        RECT 67.150 180.030 67.470 180.090 ;
        RECT 83.710 180.030 84.030 180.090 ;
        RECT 86.470 180.030 86.790 180.090 ;
        RECT 89.705 180.030 89.995 180.075 ;
        RECT 102.110 180.030 102.430 180.090 ;
        RECT 103.045 180.030 103.335 180.075 ;
        RECT 67.150 179.890 69.220 180.030 ;
        RECT 67.150 179.830 67.470 179.890 ;
        RECT 50.605 179.505 50.895 179.735 ;
        RECT 51.985 179.505 52.275 179.735 ;
        RECT 52.905 179.690 53.195 179.735 ;
        RECT 53.825 179.690 54.115 179.735 ;
        RECT 52.905 179.550 54.115 179.690 ;
        RECT 52.905 179.505 53.195 179.550 ;
        RECT 53.825 179.505 54.115 179.550 ;
        RECT 54.270 179.690 54.590 179.750 ;
        RECT 57.490 179.690 57.810 179.750 ;
        RECT 54.270 179.550 57.810 179.690 ;
        RECT 49.670 178.810 49.990 179.070 ;
        RECT 50.680 179.010 50.820 179.505 ;
        RECT 52.060 179.350 52.200 179.505 ;
        RECT 54.270 179.490 54.590 179.550 ;
        RECT 57.490 179.490 57.810 179.550 ;
        RECT 62.550 179.690 62.870 179.750 ;
        RECT 64.850 179.690 65.170 179.750 ;
        RECT 69.080 179.735 69.220 179.890 ;
        RECT 72.760 179.890 86.790 180.030 ;
        RECT 72.760 179.735 72.900 179.890 ;
        RECT 83.710 179.830 84.030 179.890 ;
        RECT 86.470 179.830 86.790 179.890 ;
        RECT 87.250 179.890 94.060 180.030 ;
        RECT 62.550 179.550 65.170 179.690 ;
        RECT 62.550 179.490 62.870 179.550 ;
        RECT 64.850 179.490 65.170 179.550 ;
        RECT 69.005 179.505 69.295 179.735 ;
        RECT 72.685 179.505 72.975 179.735 ;
        RECT 75.905 179.690 76.195 179.735 ;
        RECT 76.810 179.690 77.130 179.750 ;
        RECT 75.905 179.550 77.130 179.690 ;
        RECT 75.905 179.505 76.195 179.550 ;
        RECT 76.810 179.490 77.130 179.550 ;
        RECT 81.870 179.690 82.190 179.750 ;
        RECT 84.630 179.690 84.950 179.750 ;
        RECT 81.870 179.550 84.950 179.690 ;
        RECT 81.870 179.490 82.190 179.550 ;
        RECT 84.630 179.490 84.950 179.550 ;
        RECT 86.010 179.690 86.330 179.750 ;
        RECT 87.250 179.690 87.390 179.890 ;
        RECT 89.705 179.845 89.995 179.890 ;
        RECT 92.925 179.690 93.215 179.735 ;
        RECT 86.010 179.550 87.390 179.690 ;
        RECT 92.540 179.550 93.215 179.690 ;
        RECT 86.010 179.490 86.330 179.550 ;
        RECT 52.430 179.350 52.750 179.410 ;
        RECT 60.250 179.350 60.570 179.410 ;
        RECT 52.060 179.210 60.570 179.350 ;
        RECT 52.430 179.150 52.750 179.210 ;
        RECT 60.250 179.150 60.570 179.210 ;
        RECT 61.170 179.350 61.490 179.410 ;
        RECT 74.985 179.350 75.275 179.395 ;
        RECT 75.430 179.350 75.750 179.410 ;
        RECT 61.170 179.210 75.750 179.350 ;
        RECT 61.170 179.150 61.490 179.210 ;
        RECT 74.985 179.165 75.275 179.210 ;
        RECT 75.430 179.150 75.750 179.210 ;
        RECT 80.030 179.350 80.350 179.410 ;
        RECT 89.690 179.350 90.010 179.410 ;
        RECT 80.030 179.210 90.010 179.350 ;
        RECT 80.030 179.150 80.350 179.210 ;
        RECT 89.690 179.150 90.010 179.210 ;
        RECT 90.150 179.350 90.470 179.410 ;
        RECT 90.150 179.210 91.760 179.350 ;
        RECT 90.150 179.150 90.470 179.210 ;
        RECT 91.620 179.070 91.760 179.210 ;
        RECT 53.810 179.010 54.130 179.070 ;
        RECT 50.680 178.870 54.130 179.010 ;
        RECT 53.810 178.810 54.130 178.870 ;
        RECT 65.310 178.810 65.630 179.070 ;
        RECT 66.690 179.010 67.010 179.070 ;
        RECT 68.085 179.010 68.375 179.055 ;
        RECT 66.690 178.870 68.375 179.010 ;
        RECT 66.690 178.810 67.010 178.870 ;
        RECT 68.085 178.825 68.375 178.870 ;
        RECT 90.610 178.810 90.930 179.070 ;
        RECT 91.530 178.810 91.850 179.070 ;
        RECT 92.540 179.055 92.680 179.550 ;
        RECT 92.925 179.505 93.215 179.550 ;
        RECT 93.920 179.350 94.060 179.890 ;
        RECT 99.900 179.890 103.335 180.030 ;
        RECT 99.900 179.750 100.040 179.890 ;
        RECT 102.110 179.830 102.430 179.890 ;
        RECT 103.045 179.845 103.335 179.890 ;
        RECT 109.025 180.030 109.315 180.075 ;
        RECT 109.470 180.030 109.790 180.090 ;
        RECT 110.480 180.075 110.620 180.570 ;
        RECT 109.025 179.890 109.790 180.030 ;
        RECT 109.025 179.845 109.315 179.890 ;
        RECT 109.470 179.830 109.790 179.890 ;
        RECT 110.405 180.030 110.695 180.075 ;
        RECT 113.610 180.030 113.930 180.090 ;
        RECT 110.405 179.890 113.930 180.030 ;
        RECT 110.405 179.845 110.695 179.890 ;
        RECT 113.610 179.830 113.930 179.890 ;
        RECT 96.130 179.690 96.450 179.750 ;
        RECT 96.605 179.690 96.895 179.735 ;
        RECT 96.130 179.550 96.895 179.690 ;
        RECT 96.130 179.490 96.450 179.550 ;
        RECT 96.605 179.505 96.895 179.550 ;
        RECT 99.810 179.490 100.130 179.750 ;
        RECT 107.185 179.690 107.475 179.735 ;
        RECT 107.630 179.690 107.950 179.750 ;
        RECT 107.185 179.550 107.950 179.690 ;
        RECT 107.185 179.505 107.475 179.550 ;
        RECT 107.630 179.490 107.950 179.550 ;
        RECT 108.550 179.490 108.870 179.750 ;
        RECT 102.125 179.350 102.415 179.395 ;
        RECT 108.640 179.350 108.780 179.490 ;
        RECT 93.920 179.210 100.500 179.350 ;
        RECT 100.360 179.070 100.500 179.210 ;
        RECT 102.125 179.210 108.780 179.350 ;
        RECT 102.125 179.165 102.415 179.210 ;
        RECT 92.465 178.825 92.755 179.055 ;
        RECT 94.290 179.010 94.610 179.070 ;
        RECT 98.445 179.010 98.735 179.055 ;
        RECT 94.290 178.870 98.735 179.010 ;
        RECT 94.290 178.810 94.610 178.870 ;
        RECT 98.445 178.825 98.735 178.870 ;
        RECT 100.270 178.810 100.590 179.070 ;
        RECT 100.730 179.010 101.050 179.070 ;
        RECT 102.200 179.010 102.340 179.165 ;
        RECT 100.730 178.870 102.340 179.010 ;
        RECT 100.730 178.810 101.050 178.870 ;
        RECT 102.570 178.810 102.890 179.070 ;
        RECT 104.410 178.810 104.730 179.070 ;
        RECT 107.645 179.010 107.935 179.055 ;
        RECT 108.550 179.010 108.870 179.070 ;
        RECT 107.645 178.870 108.870 179.010 ;
        RECT 107.645 178.825 107.935 178.870 ;
        RECT 108.550 178.810 108.870 178.870 ;
        RECT 49.670 177.790 49.990 178.050 ;
        RECT 58.410 177.790 58.730 178.050 ;
        RECT 60.265 177.990 60.555 178.035 ;
        RECT 62.090 177.990 62.410 178.050 ;
        RECT 60.265 177.850 62.410 177.990 ;
        RECT 60.265 177.805 60.555 177.850 ;
        RECT 62.090 177.790 62.410 177.850 ;
        RECT 63.470 177.790 63.790 178.050 ;
        RECT 75.890 177.790 76.210 178.050 ;
        RECT 78.205 177.990 78.495 178.035 ;
        RECT 84.170 177.990 84.490 178.050 ;
        RECT 78.205 177.850 84.490 177.990 ;
        RECT 78.205 177.805 78.495 177.850 ;
        RECT 84.170 177.790 84.490 177.850 ;
        RECT 89.230 177.990 89.550 178.050 ;
        RECT 93.845 177.990 94.135 178.035 ;
        RECT 95.210 177.990 95.530 178.050 ;
        RECT 89.230 177.850 94.135 177.990 ;
        RECT 89.230 177.790 89.550 177.850 ;
        RECT 93.845 177.805 94.135 177.850 ;
        RECT 94.840 177.850 95.530 177.990 ;
        RECT 49.760 177.310 49.900 177.790 ;
        RECT 65.310 177.650 65.630 177.710 ;
        RECT 80.045 177.650 80.335 177.695 ;
        RECT 65.310 177.510 80.335 177.650 ;
        RECT 65.310 177.450 65.630 177.510 ;
        RECT 80.045 177.465 80.335 177.510 ;
        RECT 81.420 177.650 81.710 177.695 ;
        RECT 82.340 177.650 82.630 177.695 ;
        RECT 87.860 177.650 88.150 177.695 ;
        RECT 91.990 177.650 92.310 177.710 ;
        RECT 81.420 177.510 88.150 177.650 ;
        RECT 81.420 177.465 81.710 177.510 ;
        RECT 82.340 177.465 82.630 177.510 ;
        RECT 87.860 177.465 88.150 177.510 ;
        RECT 90.240 177.510 92.310 177.650 ;
        RECT 50.605 177.310 50.895 177.355 ;
        RECT 49.760 177.170 50.895 177.310 ;
        RECT 50.605 177.125 50.895 177.170 ;
        RECT 63.025 177.125 63.315 177.355 ;
        RECT 69.005 177.125 69.295 177.355 ;
        RECT 51.510 176.770 51.830 177.030 ;
        RECT 51.985 176.970 52.275 177.015 ;
        RECT 57.490 176.970 57.810 177.030 ;
        RECT 51.985 176.830 57.810 176.970 ;
        RECT 51.985 176.785 52.275 176.830 ;
        RECT 57.490 176.770 57.810 176.830 ;
        RECT 60.710 176.770 61.030 177.030 ;
        RECT 61.170 176.970 61.490 177.030 ;
        RECT 63.100 176.970 63.240 177.125 ;
        RECT 66.230 176.970 66.550 177.030 ;
        RECT 68.085 176.970 68.375 177.015 ;
        RECT 61.170 176.830 68.375 176.970 ;
        RECT 69.080 176.970 69.220 177.125 ;
        RECT 73.130 177.110 73.450 177.370 ;
        RECT 84.170 177.355 84.490 177.370 ;
        RECT 77.745 177.310 78.035 177.355 ;
        RECT 80.915 177.310 81.205 177.355 ;
        RECT 82.755 177.310 83.045 177.355 ;
        RECT 77.745 177.170 80.720 177.310 ;
        RECT 77.745 177.125 78.035 177.170 ;
        RECT 73.220 176.970 73.360 177.110 ;
        RECT 78.665 176.970 78.955 177.015 ;
        RECT 80.030 176.970 80.350 177.030 ;
        RECT 69.080 176.830 73.360 176.970 ;
        RECT 78.280 176.830 80.350 176.970 ;
        RECT 61.170 176.770 61.490 176.830 ;
        RECT 66.230 176.770 66.550 176.830 ;
        RECT 68.085 176.785 68.375 176.830 ;
        RECT 49.685 176.630 49.975 176.675 ;
        RECT 56.570 176.630 56.890 176.690 ;
        RECT 49.685 176.490 56.890 176.630 ;
        RECT 49.685 176.445 49.975 176.490 ;
        RECT 56.570 176.430 56.890 176.490 ;
        RECT 63.470 176.290 63.790 176.350 ;
        RECT 74.050 176.290 74.370 176.350 ;
        RECT 78.280 176.290 78.420 176.830 ;
        RECT 78.665 176.785 78.955 176.830 ;
        RECT 80.030 176.770 80.350 176.830 ;
        RECT 63.470 176.150 78.420 176.290 ;
        RECT 80.580 176.290 80.720 177.170 ;
        RECT 80.915 177.170 83.045 177.310 ;
        RECT 80.915 177.125 81.205 177.170 ;
        RECT 82.755 177.125 83.045 177.170 ;
        RECT 84.060 177.125 84.490 177.355 ;
        RECT 84.170 177.110 84.490 177.125 ;
        RECT 84.630 177.110 84.950 177.370 ;
        RECT 85.100 177.310 85.390 177.355 ;
        RECT 86.940 177.310 87.230 177.355 ;
        RECT 85.100 177.170 87.230 177.310 ;
        RECT 85.100 177.125 85.390 177.170 ;
        RECT 86.940 177.125 87.230 177.170 ;
        RECT 88.325 177.310 88.615 177.355 ;
        RECT 89.705 177.310 89.995 177.355 ;
        RECT 88.325 177.170 89.995 177.310 ;
        RECT 88.325 177.125 88.615 177.170 ;
        RECT 89.705 177.125 89.995 177.170 ;
        RECT 82.330 176.970 82.650 177.030 ;
        RECT 83.265 176.970 83.555 177.015 ;
        RECT 82.330 176.830 83.555 176.970 ;
        RECT 82.330 176.770 82.650 176.830 ;
        RECT 83.265 176.785 83.555 176.830 ;
        RECT 86.025 176.970 86.315 177.015 ;
        RECT 88.770 176.970 89.090 177.030 ;
        RECT 86.025 176.830 89.090 176.970 ;
        RECT 86.025 176.785 86.315 176.830 ;
        RECT 88.770 176.770 89.090 176.830 ;
        RECT 89.245 176.970 89.535 177.015 ;
        RECT 90.240 176.970 90.380 177.510 ;
        RECT 91.990 177.450 92.310 177.510 ;
        RECT 90.625 177.310 90.915 177.355 ;
        RECT 94.840 177.310 94.980 177.850 ;
        RECT 95.210 177.790 95.530 177.850 ;
        RECT 96.590 177.990 96.910 178.050 ;
        RECT 108.105 177.990 108.395 178.035 ;
        RECT 109.930 177.990 110.250 178.050 ;
        RECT 96.590 177.850 110.250 177.990 ;
        RECT 96.590 177.790 96.910 177.850 ;
        RECT 108.105 177.805 108.395 177.850 ;
        RECT 109.930 177.790 110.250 177.850 ;
        RECT 96.130 177.650 96.450 177.710 ;
        RECT 99.350 177.650 99.670 177.710 ;
        RECT 105.345 177.650 105.635 177.695 ;
        RECT 96.130 177.510 98.660 177.650 ;
        RECT 96.130 177.450 96.450 177.510 ;
        RECT 90.625 177.170 94.980 177.310 ;
        RECT 95.210 177.310 95.530 177.370 ;
        RECT 98.520 177.355 98.660 177.510 ;
        RECT 99.350 177.510 105.635 177.650 ;
        RECT 99.350 177.450 99.670 177.510 ;
        RECT 105.345 177.465 105.635 177.510 ;
        RECT 95.685 177.310 95.975 177.355 ;
        RECT 95.210 177.170 95.975 177.310 ;
        RECT 90.625 177.125 90.915 177.170 ;
        RECT 95.210 177.110 95.530 177.170 ;
        RECT 95.685 177.125 95.975 177.170 ;
        RECT 98.445 177.310 98.735 177.355 ;
        RECT 102.110 177.310 102.430 177.370 ;
        RECT 98.445 177.170 102.430 177.310 ;
        RECT 98.445 177.125 98.735 177.170 ;
        RECT 102.110 177.110 102.430 177.170 ;
        RECT 103.490 177.110 103.810 177.370 ;
        RECT 104.870 177.110 105.190 177.370 ;
        RECT 112.230 177.310 112.550 177.370 ;
        RECT 113.625 177.310 113.915 177.355 ;
        RECT 112.230 177.170 113.915 177.310 ;
        RECT 112.230 177.110 112.550 177.170 ;
        RECT 113.625 177.125 113.915 177.170 ;
        RECT 89.245 176.830 90.380 176.970 ;
        RECT 96.145 176.970 96.435 177.015 ;
        RECT 96.590 176.970 96.910 177.030 ;
        RECT 96.145 176.830 96.910 176.970 ;
        RECT 89.245 176.785 89.535 176.830 ;
        RECT 96.145 176.785 96.435 176.830 ;
        RECT 96.590 176.770 96.910 176.830 ;
        RECT 97.065 176.970 97.355 177.015 ;
        RECT 99.810 176.970 100.130 177.030 ;
        RECT 97.065 176.830 100.130 176.970 ;
        RECT 97.065 176.785 97.355 176.830 ;
        RECT 99.810 176.770 100.130 176.830 ;
        RECT 100.270 176.970 100.590 177.030 ;
        RECT 101.205 176.970 101.495 177.015 ;
        RECT 103.580 176.970 103.720 177.110 ;
        RECT 100.270 176.830 103.720 176.970 ;
        RECT 100.270 176.770 100.590 176.830 ;
        RECT 101.205 176.785 101.495 176.830 ;
        RECT 104.410 176.770 104.730 177.030 ;
        RECT 105.805 176.785 106.095 177.015 ;
        RECT 81.835 176.630 82.125 176.675 ;
        RECT 85.065 176.630 85.355 176.675 ;
        RECT 81.835 176.490 85.355 176.630 ;
        RECT 81.835 176.445 82.125 176.490 ;
        RECT 85.065 176.445 85.355 176.490 ;
        RECT 92.910 176.630 93.230 176.690 ;
        RECT 104.500 176.630 104.640 176.770 ;
        RECT 92.910 176.490 104.640 176.630 ;
        RECT 92.910 176.430 93.230 176.490 ;
        RECT 89.230 176.290 89.550 176.350 ;
        RECT 80.580 176.150 89.550 176.290 ;
        RECT 63.470 176.090 63.790 176.150 ;
        RECT 74.050 176.090 74.370 176.150 ;
        RECT 89.230 176.090 89.550 176.150 ;
        RECT 93.370 176.290 93.690 176.350 ;
        RECT 99.350 176.290 99.670 176.350 ;
        RECT 93.370 176.150 99.670 176.290 ;
        RECT 93.370 176.090 93.690 176.150 ;
        RECT 99.350 176.090 99.670 176.150 ;
        RECT 103.030 176.090 103.350 176.350 ;
        RECT 104.410 176.290 104.730 176.350 ;
        RECT 105.880 176.290 106.020 176.785 ;
        RECT 111.310 176.770 111.630 177.030 ;
        RECT 104.410 176.150 106.020 176.290 ;
        RECT 104.410 176.090 104.730 176.150 ;
        RECT 57.505 175.270 57.795 175.315 ;
        RECT 60.710 175.270 61.030 175.330 ;
        RECT 86.010 175.270 86.330 175.330 ;
        RECT 89.690 175.270 90.010 175.330 ;
        RECT 57.505 175.130 61.030 175.270 ;
        RECT 57.505 175.085 57.795 175.130 ;
        RECT 60.710 175.070 61.030 175.130 ;
        RECT 81.960 175.130 90.010 175.270 ;
        RECT 51.525 174.930 51.815 174.975 ;
        RECT 72.670 174.930 72.990 174.990 ;
        RECT 73.605 174.930 73.895 174.975 ;
        RECT 74.050 174.930 74.370 174.990 ;
        RECT 51.525 174.790 55.880 174.930 ;
        RECT 51.525 174.745 51.815 174.790 ;
        RECT 50.145 174.590 50.435 174.635 ;
        RECT 52.430 174.590 52.750 174.650 ;
        RECT 55.740 174.635 55.880 174.790 ;
        RECT 69.080 174.790 74.370 174.930 ;
        RECT 50.145 174.450 52.750 174.590 ;
        RECT 50.145 174.405 50.435 174.450 ;
        RECT 52.430 174.390 52.750 174.450 ;
        RECT 55.665 174.405 55.955 174.635 ;
        RECT 61.170 174.590 61.490 174.650 ;
        RECT 69.080 174.635 69.220 174.790 ;
        RECT 72.670 174.730 72.990 174.790 ;
        RECT 73.605 174.745 73.895 174.790 ;
        RECT 74.050 174.730 74.370 174.790 ;
        RECT 74.565 174.930 74.855 174.975 ;
        RECT 77.795 174.930 78.085 174.975 ;
        RECT 74.565 174.790 78.085 174.930 ;
        RECT 74.565 174.745 74.855 174.790 ;
        RECT 77.795 174.745 78.085 174.790 ;
        RECT 81.960 174.635 82.100 175.130 ;
        RECT 86.010 175.070 86.330 175.130 ;
        RECT 89.690 175.070 90.010 175.130 ;
        RECT 92.005 175.270 92.295 175.315 ;
        RECT 93.370 175.270 93.690 175.330 ;
        RECT 92.005 175.130 93.690 175.270 ;
        RECT 92.005 175.085 92.295 175.130 ;
        RECT 93.370 175.070 93.690 175.130 ;
        RECT 96.590 175.270 96.910 175.330 ;
        RECT 97.525 175.270 97.815 175.315 ;
        RECT 96.590 175.130 97.815 175.270 ;
        RECT 96.590 175.070 96.910 175.130 ;
        RECT 97.525 175.085 97.815 175.130 ;
        RECT 84.630 174.730 84.950 174.990 ;
        RECT 100.360 174.790 104.180 174.930 ;
        RECT 62.565 174.590 62.855 174.635 ;
        RECT 61.170 174.450 62.855 174.590 ;
        RECT 61.170 174.390 61.490 174.450 ;
        RECT 62.565 174.405 62.855 174.450 ;
        RECT 69.005 174.405 69.295 174.635 ;
        RECT 71.075 174.590 71.365 174.635 ;
        RECT 75.570 174.590 75.860 174.635 ;
        RECT 69.540 174.450 71.365 174.590 ;
        RECT 49.685 174.250 49.975 174.295 ;
        RECT 51.970 174.250 52.290 174.310 ;
        RECT 49.685 174.110 52.290 174.250 ;
        RECT 49.685 174.065 49.975 174.110 ;
        RECT 51.970 174.050 52.290 174.110 ;
        RECT 55.190 174.250 55.510 174.310 ;
        RECT 56.125 174.250 56.415 174.295 ;
        RECT 58.870 174.250 59.190 174.310 ;
        RECT 55.190 174.110 59.190 174.250 ;
        RECT 55.190 174.050 55.510 174.110 ;
        RECT 56.125 174.065 56.415 174.110 ;
        RECT 58.870 174.050 59.190 174.110 ;
        RECT 59.330 174.050 59.650 174.310 ;
        RECT 67.610 174.250 67.930 174.310 ;
        RECT 69.540 174.250 69.680 174.450 ;
        RECT 71.075 174.405 71.365 174.450 ;
        RECT 72.300 174.450 75.860 174.590 ;
        RECT 72.300 174.310 72.440 174.450 ;
        RECT 75.570 174.405 75.860 174.450 ;
        RECT 81.885 174.405 82.175 174.635 ;
        RECT 82.345 174.590 82.635 174.635 ;
        RECT 82.790 174.590 83.110 174.650 ;
        RECT 89.230 174.590 89.550 174.650 ;
        RECT 93.385 174.590 93.675 174.635 ;
        RECT 99.810 174.590 100.130 174.650 ;
        RECT 82.345 174.450 83.110 174.590 ;
        RECT 82.345 174.405 82.635 174.450 ;
        RECT 82.790 174.390 83.110 174.450 ;
        RECT 83.800 174.450 87.390 174.590 ;
        RECT 64.020 174.110 69.680 174.250 ;
        RECT 69.910 174.250 70.230 174.310 ;
        RECT 70.385 174.250 70.675 174.295 ;
        RECT 69.910 174.110 70.675 174.250 ;
        RECT 64.020 173.955 64.160 174.110 ;
        RECT 67.610 174.050 67.930 174.110 ;
        RECT 69.910 174.050 70.230 174.110 ;
        RECT 70.385 174.065 70.675 174.110 ;
        RECT 72.210 174.050 72.530 174.310 ;
        RECT 72.690 174.250 72.980 174.295 ;
        RECT 74.530 174.250 74.820 174.295 ;
        RECT 72.690 174.110 74.820 174.250 ;
        RECT 72.690 174.065 72.980 174.110 ;
        RECT 74.530 174.065 74.820 174.110 ;
        RECT 74.970 174.050 75.290 174.310 ;
        RECT 76.350 174.050 76.670 174.310 ;
        RECT 76.875 174.250 77.165 174.295 ;
        RECT 78.715 174.250 79.005 174.295 ;
        RECT 76.875 174.110 79.005 174.250 ;
        RECT 76.875 174.065 77.165 174.110 ;
        RECT 78.715 174.065 79.005 174.110 ;
        RECT 79.585 174.250 79.875 174.295 ;
        RECT 83.800 174.250 83.940 174.450 ;
        RECT 79.585 174.110 83.940 174.250 ;
        RECT 84.630 174.250 84.950 174.310 ;
        RECT 86.025 174.250 86.315 174.295 ;
        RECT 84.630 174.110 86.315 174.250 ;
        RECT 87.250 174.250 87.390 174.450 ;
        RECT 89.230 174.450 100.130 174.590 ;
        RECT 89.230 174.390 89.550 174.450 ;
        RECT 93.385 174.405 93.675 174.450 ;
        RECT 99.810 174.390 100.130 174.450 ;
        RECT 89.705 174.250 89.995 174.295 ;
        RECT 87.250 174.110 89.995 174.250 ;
        RECT 79.585 174.065 79.875 174.110 ;
        RECT 84.630 174.050 84.950 174.110 ;
        RECT 86.025 174.065 86.315 174.110 ;
        RECT 89.705 174.065 89.995 174.110 ;
        RECT 90.150 174.050 90.470 174.310 ;
        RECT 94.290 174.050 94.610 174.310 ;
        RECT 100.360 174.250 100.500 174.790 ;
        RECT 100.745 174.590 101.035 174.635 ;
        RECT 101.650 174.590 101.970 174.650 ;
        RECT 102.570 174.590 102.890 174.650 ;
        RECT 100.745 174.450 102.890 174.590 ;
        RECT 100.745 174.405 101.035 174.450 ;
        RECT 101.650 174.390 101.970 174.450 ;
        RECT 102.570 174.390 102.890 174.450 ;
        RECT 103.030 174.390 103.350 174.650 ;
        RECT 104.040 174.635 104.180 174.790 ;
        RECT 103.965 174.405 104.255 174.635 ;
        RECT 104.410 174.390 104.730 174.650 ;
        RECT 109.470 174.590 109.790 174.650 ;
        RECT 104.960 174.450 109.790 174.590 ;
        RECT 96.220 174.110 100.500 174.250 ;
        RECT 103.120 174.250 103.260 174.390 ;
        RECT 103.505 174.250 103.795 174.295 ;
        RECT 103.120 174.110 103.795 174.250 ;
        RECT 63.945 173.910 64.235 173.955 ;
        RECT 56.200 173.770 64.235 173.910 ;
        RECT 56.200 173.630 56.340 173.770 ;
        RECT 63.945 173.725 64.235 173.770 ;
        RECT 71.770 173.910 72.060 173.955 ;
        RECT 77.290 173.910 77.580 173.955 ;
        RECT 78.210 173.910 78.500 173.955 ;
        RECT 82.805 173.910 83.095 173.955 ;
        RECT 94.380 173.910 94.520 174.050 ;
        RECT 71.770 173.770 78.500 173.910 ;
        RECT 71.770 173.725 72.060 173.770 ;
        RECT 77.290 173.725 77.580 173.770 ;
        RECT 78.210 173.725 78.500 173.770 ;
        RECT 78.740 173.770 83.095 173.910 ;
        RECT 56.110 173.370 56.430 173.630 ;
        RECT 58.410 173.370 58.730 173.630 ;
        RECT 63.470 173.370 63.790 173.630 ;
        RECT 65.770 173.370 66.090 173.630 ;
        RECT 66.230 173.370 66.550 173.630 ;
        RECT 68.070 173.370 68.390 173.630 ;
        RECT 68.545 173.570 68.835 173.615 ;
        RECT 74.970 173.570 75.290 173.630 ;
        RECT 68.545 173.430 75.290 173.570 ;
        RECT 68.545 173.385 68.835 173.430 ;
        RECT 74.970 173.370 75.290 173.430 ;
        RECT 76.350 173.570 76.670 173.630 ;
        RECT 78.740 173.570 78.880 173.770 ;
        RECT 82.805 173.725 83.095 173.770 ;
        RECT 87.250 173.770 94.520 173.910 ;
        RECT 76.350 173.430 78.880 173.570 ;
        RECT 76.350 173.370 76.670 173.430 ;
        RECT 85.090 173.370 85.410 173.630 ;
        RECT 86.010 173.570 86.330 173.630 ;
        RECT 87.250 173.570 87.390 173.770 ;
        RECT 86.010 173.430 87.390 173.570 ;
        RECT 87.850 173.570 88.170 173.630 ;
        RECT 93.830 173.570 94.150 173.630 ;
        RECT 87.850 173.430 94.150 173.570 ;
        RECT 86.010 173.370 86.330 173.430 ;
        RECT 87.850 173.370 88.170 173.430 ;
        RECT 93.830 173.370 94.150 173.430 ;
        RECT 94.290 173.370 94.610 173.630 ;
        RECT 96.220 173.615 96.360 174.110 ;
        RECT 103.505 174.065 103.795 174.110 ;
        RECT 98.430 173.910 98.750 173.970 ;
        RECT 99.365 173.910 99.655 173.955 ;
        RECT 104.960 173.910 105.100 174.450 ;
        RECT 109.470 174.390 109.790 174.450 ;
        RECT 112.230 174.590 112.550 174.650 ;
        RECT 112.705 174.590 112.995 174.635 ;
        RECT 112.230 174.450 112.995 174.590 ;
        RECT 112.230 174.390 112.550 174.450 ;
        RECT 112.705 174.405 112.995 174.450 ;
        RECT 108.550 174.050 108.870 174.310 ;
        RECT 109.010 174.050 109.330 174.310 ;
        RECT 98.430 173.770 105.100 173.910 ;
        RECT 105.790 173.910 106.110 173.970 ;
        RECT 109.100 173.910 109.240 174.050 ;
        RECT 105.790 173.770 108.780 173.910 ;
        RECT 109.100 173.770 112.000 173.910 ;
        RECT 98.430 173.710 98.750 173.770 ;
        RECT 99.365 173.725 99.655 173.770 ;
        RECT 105.790 173.710 106.110 173.770 ;
        RECT 96.145 173.385 96.435 173.615 ;
        RECT 99.810 173.370 100.130 173.630 ;
        RECT 100.270 173.570 100.590 173.630 ;
        RECT 101.665 173.570 101.955 173.615 ;
        RECT 100.270 173.430 101.955 173.570 ;
        RECT 100.270 173.370 100.590 173.430 ;
        RECT 101.665 173.385 101.955 173.430 ;
        RECT 104.870 173.570 105.190 173.630 ;
        RECT 106.725 173.570 107.015 173.615 ;
        RECT 104.870 173.430 107.015 173.570 ;
        RECT 108.640 173.570 108.780 173.770 ;
        RECT 111.860 173.630 112.000 173.770 ;
        RECT 109.025 173.570 109.315 173.615 ;
        RECT 108.640 173.430 109.315 173.570 ;
        RECT 104.870 173.370 105.190 173.430 ;
        RECT 106.725 173.385 107.015 173.430 ;
        RECT 109.025 173.385 109.315 173.430 ;
        RECT 111.770 173.370 112.090 173.630 ;
        RECT 113.150 173.570 113.470 173.630 ;
        RECT 114.530 173.570 114.850 173.630 ;
        RECT 113.150 173.430 114.850 173.570 ;
        RECT 113.150 173.370 113.470 173.430 ;
        RECT 114.530 173.370 114.850 173.430 ;
        RECT 56.125 172.550 56.415 172.595 ;
        RECT 57.030 172.550 57.350 172.610 ;
        RECT 68.070 172.550 68.390 172.610 ;
        RECT 72.210 172.550 72.530 172.610 ;
        RECT 56.125 172.410 57.350 172.550 ;
        RECT 56.125 172.365 56.415 172.410 ;
        RECT 57.030 172.350 57.350 172.410 ;
        RECT 58.040 172.410 72.530 172.550 ;
        RECT 44.610 171.870 44.930 171.930 ;
        RECT 58.040 171.915 58.180 172.410 ;
        RECT 68.070 172.350 68.390 172.410 ;
        RECT 72.210 172.350 72.530 172.410 ;
        RECT 83.250 172.350 83.570 172.610 ;
        RECT 88.310 172.350 88.630 172.610 ;
        RECT 89.230 172.550 89.550 172.610 ;
        RECT 90.165 172.550 90.455 172.595 ;
        RECT 89.230 172.410 90.455 172.550 ;
        RECT 89.230 172.350 89.550 172.410 ;
        RECT 90.165 172.365 90.455 172.410 ;
        RECT 94.750 172.550 95.070 172.610 ;
        RECT 97.970 172.550 98.290 172.610 ;
        RECT 94.750 172.410 98.290 172.550 ;
        RECT 94.750 172.350 95.070 172.410 ;
        RECT 97.970 172.350 98.290 172.410 ;
        RECT 103.950 172.550 104.270 172.610 ;
        RECT 108.550 172.550 108.870 172.610 ;
        RECT 114.085 172.550 114.375 172.595 ;
        RECT 103.950 172.410 106.020 172.550 ;
        RECT 103.950 172.350 104.270 172.410 ;
        RECT 64.390 172.210 64.710 172.270 ;
        RECT 69.910 172.210 70.230 172.270 ;
        RECT 72.670 172.210 72.990 172.270 ;
        RECT 64.390 172.070 68.760 172.210 ;
        RECT 64.390 172.010 64.710 172.070 ;
        RECT 57.965 171.870 58.255 171.915 ;
        RECT 44.610 171.730 58.255 171.870 ;
        RECT 44.610 171.670 44.930 171.730 ;
        RECT 57.965 171.685 58.255 171.730 ;
        RECT 58.870 171.870 59.190 171.930 ;
        RECT 63.945 171.870 64.235 171.915 ;
        RECT 58.870 171.730 64.235 171.870 ;
        RECT 58.870 171.670 59.190 171.730 ;
        RECT 63.945 171.685 64.235 171.730 ;
        RECT 64.865 171.870 65.155 171.915 ;
        RECT 65.770 171.870 66.090 171.930 ;
        RECT 64.865 171.730 66.090 171.870 ;
        RECT 64.865 171.685 65.155 171.730 ;
        RECT 54.270 171.530 54.590 171.590 ;
        RECT 58.425 171.530 58.715 171.575 ;
        RECT 54.270 171.390 58.715 171.530 ;
        RECT 54.270 171.330 54.590 171.390 ;
        RECT 58.425 171.345 58.715 171.390 ;
        RECT 59.345 171.530 59.635 171.575 ;
        RECT 60.710 171.530 61.030 171.590 ;
        RECT 59.345 171.390 61.030 171.530 ;
        RECT 64.020 171.530 64.160 171.685 ;
        RECT 65.770 171.670 66.090 171.730 ;
        RECT 66.230 171.870 66.550 171.930 ;
        RECT 68.085 171.870 68.375 171.915 ;
        RECT 66.230 171.730 68.375 171.870 ;
        RECT 68.620 171.870 68.760 172.070 ;
        RECT 69.910 172.070 72.990 172.210 ;
        RECT 69.910 172.010 70.230 172.070 ;
        RECT 72.670 172.010 72.990 172.070 ;
        RECT 75.890 172.210 76.210 172.270 ;
        RECT 87.390 172.210 87.710 172.270 ;
        RECT 88.400 172.210 88.540 172.350 ;
        RECT 75.890 172.070 87.710 172.210 ;
        RECT 75.890 172.010 76.210 172.070 ;
        RECT 87.390 172.010 87.710 172.070 ;
        RECT 87.940 172.070 88.540 172.210 ;
        RECT 101.650 172.210 101.970 172.270 ;
        RECT 104.410 172.210 104.730 172.270 ;
        RECT 101.650 172.070 104.730 172.210 ;
        RECT 82.790 171.870 83.110 171.930 ;
        RECT 68.620 171.730 83.110 171.870 ;
        RECT 66.230 171.670 66.550 171.730 ;
        RECT 68.085 171.685 68.375 171.730 ;
        RECT 82.790 171.670 83.110 171.730 ;
        RECT 86.930 171.670 87.250 171.930 ;
        RECT 87.940 171.915 88.080 172.070 ;
        RECT 101.650 172.010 101.970 172.070 ;
        RECT 104.410 172.010 104.730 172.070 ;
        RECT 87.865 171.685 88.155 171.915 ;
        RECT 97.985 171.870 98.275 171.915 ;
        RECT 98.430 171.870 98.750 171.930 ;
        RECT 97.985 171.730 98.750 171.870 ;
        RECT 97.985 171.685 98.275 171.730 ;
        RECT 98.430 171.670 98.750 171.730 ;
        RECT 98.890 171.670 99.210 171.930 ;
        RECT 104.870 171.670 105.190 171.930 ;
        RECT 105.880 171.915 106.020 172.410 ;
        RECT 108.550 172.410 114.375 172.550 ;
        RECT 108.550 172.350 108.870 172.410 ;
        RECT 114.085 172.365 114.375 172.410 ;
        RECT 106.270 172.210 106.560 172.255 ;
        RECT 111.790 172.210 112.080 172.255 ;
        RECT 112.710 172.210 113.000 172.255 ;
        RECT 106.270 172.070 113.000 172.210 ;
        RECT 106.270 172.025 106.560 172.070 ;
        RECT 111.790 172.025 112.080 172.070 ;
        RECT 112.710 172.025 113.000 172.070 ;
        RECT 105.805 171.685 106.095 171.915 ;
        RECT 107.190 171.870 107.480 171.915 ;
        RECT 109.030 171.870 109.320 171.915 ;
        RECT 107.190 171.730 109.320 171.870 ;
        RECT 107.190 171.685 107.480 171.730 ;
        RECT 109.030 171.685 109.320 171.730 ;
        RECT 109.470 171.670 109.790 171.930 ;
        RECT 111.375 171.870 111.665 171.915 ;
        RECT 113.215 171.870 113.505 171.915 ;
        RECT 111.375 171.730 113.505 171.870 ;
        RECT 111.375 171.685 111.665 171.730 ;
        RECT 113.215 171.685 113.505 171.730 ;
        RECT 66.690 171.530 67.010 171.590 ;
        RECT 64.020 171.390 67.010 171.530 ;
        RECT 59.345 171.345 59.635 171.390 ;
        RECT 60.710 171.330 61.030 171.390 ;
        RECT 66.690 171.330 67.010 171.390 ;
        RECT 84.185 171.530 84.475 171.575 ;
        RECT 95.210 171.530 95.530 171.590 ;
        RECT 110.070 171.530 110.360 171.575 ;
        RECT 84.185 171.390 88.540 171.530 ;
        RECT 84.185 171.345 84.475 171.390 ;
        RECT 65.785 171.190 66.075 171.235 ;
        RECT 87.850 171.190 88.170 171.250 ;
        RECT 65.785 171.050 88.170 171.190 ;
        RECT 88.400 171.190 88.540 171.390 ;
        RECT 95.210 171.390 110.360 171.530 ;
        RECT 95.210 171.330 95.530 171.390 ;
        RECT 110.070 171.345 110.360 171.390 ;
        RECT 110.865 171.530 111.155 171.575 ;
        RECT 110.865 171.390 112.920 171.530 ;
        RECT 110.865 171.345 111.155 171.390 ;
        RECT 94.750 171.190 95.070 171.250 ;
        RECT 88.400 171.050 95.070 171.190 ;
        RECT 65.785 171.005 66.075 171.050 ;
        RECT 87.850 170.990 88.170 171.050 ;
        RECT 94.750 170.990 95.070 171.050 ;
        RECT 99.810 170.990 100.130 171.250 ;
        RECT 100.270 171.190 100.590 171.250 ;
        RECT 108.105 171.190 108.395 171.235 ;
        RECT 100.270 171.050 108.395 171.190 ;
        RECT 100.270 170.990 100.590 171.050 ;
        RECT 108.105 171.005 108.395 171.050 ;
        RECT 109.065 171.190 109.355 171.235 ;
        RECT 112.295 171.190 112.585 171.235 ;
        RECT 109.065 171.050 112.585 171.190 ;
        RECT 109.065 171.005 109.355 171.050 ;
        RECT 112.295 171.005 112.585 171.050 ;
        RECT 54.730 170.850 55.050 170.910 ;
        RECT 63.025 170.850 63.315 170.895 ;
        RECT 54.730 170.710 63.315 170.850 ;
        RECT 54.730 170.650 55.050 170.710 ;
        RECT 63.025 170.665 63.315 170.710 ;
        RECT 68.070 170.850 68.390 170.910 ;
        RECT 69.005 170.850 69.295 170.895 ;
        RECT 68.070 170.710 69.295 170.850 ;
        RECT 68.070 170.650 68.390 170.710 ;
        RECT 69.005 170.665 69.295 170.710 ;
        RECT 80.950 170.650 81.270 170.910 ;
        RECT 81.410 170.850 81.730 170.910 ;
        RECT 87.390 170.850 87.710 170.910 ;
        RECT 81.410 170.710 87.710 170.850 ;
        RECT 81.410 170.650 81.730 170.710 ;
        RECT 87.390 170.650 87.710 170.710 ;
        RECT 88.325 170.850 88.615 170.895 ;
        RECT 93.830 170.850 94.150 170.910 ;
        RECT 88.325 170.710 94.150 170.850 ;
        RECT 88.325 170.665 88.615 170.710 ;
        RECT 93.830 170.650 94.150 170.710 ;
        RECT 99.365 170.850 99.655 170.895 ;
        RECT 99.900 170.850 100.040 170.990 ;
        RECT 99.365 170.710 100.040 170.850 ;
        RECT 104.870 170.850 105.190 170.910 ;
        RECT 105.790 170.850 106.110 170.910 ;
        RECT 104.870 170.710 106.110 170.850 ;
        RECT 99.365 170.665 99.655 170.710 ;
        RECT 104.870 170.650 105.190 170.710 ;
        RECT 105.790 170.650 106.110 170.710 ;
        RECT 109.930 170.850 110.250 170.910 ;
        RECT 112.780 170.850 112.920 171.390 ;
        RECT 109.930 170.710 112.920 170.850 ;
        RECT 109.930 170.650 110.250 170.710 ;
        RECT 63.930 169.630 64.250 169.890 ;
        RECT 70.845 169.830 71.135 169.875 ;
        RECT 75.890 169.830 76.210 169.890 ;
        RECT 70.845 169.690 76.210 169.830 ;
        RECT 70.845 169.645 71.135 169.690 ;
        RECT 75.890 169.630 76.210 169.690 ;
        RECT 83.250 169.830 83.570 169.890 ;
        RECT 90.150 169.830 90.470 169.890 ;
        RECT 91.085 169.830 91.375 169.875 ;
        RECT 83.250 169.690 85.780 169.830 ;
        RECT 83.250 169.630 83.570 169.690 ;
        RECT 74.050 169.490 74.370 169.550 ;
        RECT 74.050 169.350 74.740 169.490 ;
        RECT 74.050 169.290 74.370 169.350 ;
        RECT 60.710 168.950 61.030 169.210 ;
        RECT 67.610 169.150 67.930 169.210 ;
        RECT 72.670 169.150 72.990 169.210 ;
        RECT 74.600 169.195 74.740 169.350 ;
        RECT 67.610 169.010 70.140 169.150 ;
        RECT 67.610 168.950 67.930 169.010 ;
        RECT 55.190 168.810 55.510 168.870 ;
        RECT 68.070 168.810 68.390 168.870 ;
        RECT 55.190 168.670 68.390 168.810 ;
        RECT 55.190 168.610 55.510 168.670 ;
        RECT 68.070 168.610 68.390 168.670 ;
        RECT 68.530 168.610 68.850 168.870 ;
        RECT 69.465 168.625 69.755 168.855 ;
        RECT 70.000 168.810 70.140 169.010 ;
        RECT 72.670 169.010 74.280 169.150 ;
        RECT 72.670 168.950 72.990 169.010 ;
        RECT 74.140 168.855 74.280 169.010 ;
        RECT 74.525 168.965 74.815 169.195 ;
        RECT 81.410 168.950 81.730 169.210 ;
        RECT 83.710 169.150 84.030 169.210 ;
        RECT 85.105 169.150 85.395 169.195 ;
        RECT 83.710 169.010 85.395 169.150 ;
        RECT 85.640 169.150 85.780 169.690 ;
        RECT 90.150 169.690 91.375 169.830 ;
        RECT 90.150 169.630 90.470 169.690 ;
        RECT 91.085 169.645 91.375 169.690 ;
        RECT 95.685 169.830 95.975 169.875 ;
        RECT 98.890 169.830 99.210 169.890 ;
        RECT 95.685 169.690 99.210 169.830 ;
        RECT 95.685 169.645 95.975 169.690 ;
        RECT 98.890 169.630 99.210 169.690 ;
        RECT 103.490 169.830 103.810 169.890 ;
        RECT 106.725 169.830 107.015 169.875 ;
        RECT 103.490 169.690 107.015 169.830 ;
        RECT 103.490 169.630 103.810 169.690 ;
        RECT 106.725 169.645 107.015 169.690 ;
        RECT 86.065 169.490 86.355 169.535 ;
        RECT 89.295 169.490 89.585 169.535 ;
        RECT 94.290 169.490 94.610 169.550 ;
        RECT 86.065 169.350 89.585 169.490 ;
        RECT 86.065 169.305 86.355 169.350 ;
        RECT 89.295 169.305 89.585 169.350 ;
        RECT 93.000 169.350 94.610 169.490 ;
        RECT 86.930 169.195 87.250 169.210 ;
        RECT 93.000 169.195 93.140 169.350 ;
        RECT 94.290 169.290 94.610 169.350 ;
        RECT 100.785 169.490 101.075 169.535 ;
        RECT 104.015 169.490 104.305 169.535 ;
        RECT 100.785 169.350 104.305 169.490 ;
        RECT 100.785 169.305 101.075 169.350 ;
        RECT 104.015 169.305 104.305 169.350 ;
        RECT 104.870 169.490 105.190 169.550 ;
        RECT 105.805 169.490 106.095 169.535 ;
        RECT 110.865 169.490 111.155 169.535 ;
        RECT 104.870 169.350 106.095 169.490 ;
        RECT 104.870 169.290 105.190 169.350 ;
        RECT 105.805 169.305 106.095 169.350 ;
        RECT 109.100 169.350 111.155 169.490 ;
        RECT 85.640 169.010 86.700 169.150 ;
        RECT 83.710 168.950 84.030 169.010 ;
        RECT 85.105 168.965 85.395 169.010 ;
        RECT 73.605 168.810 73.895 168.855 ;
        RECT 70.000 168.670 73.895 168.810 ;
        RECT 73.605 168.625 73.895 168.670 ;
        RECT 74.065 168.810 74.355 168.855 ;
        RECT 81.500 168.810 81.640 168.950 ;
        RECT 74.065 168.670 81.640 168.810 ;
        RECT 74.065 168.625 74.355 168.670 ;
        RECT 81.885 168.625 82.175 168.855 ;
        RECT 64.390 168.470 64.710 168.530 ;
        RECT 62.180 168.330 64.710 168.470 ;
        RECT 69.540 168.470 69.680 168.625 ;
        RECT 76.810 168.470 77.130 168.530 ;
        RECT 81.410 168.470 81.730 168.530 ;
        RECT 69.540 168.330 81.730 168.470 ;
        RECT 57.950 168.130 58.270 168.190 ;
        RECT 62.180 168.175 62.320 168.330 ;
        RECT 64.390 168.270 64.710 168.330 ;
        RECT 76.810 168.270 77.130 168.330 ;
        RECT 81.410 168.270 81.730 168.330 ;
        RECT 61.645 168.130 61.935 168.175 ;
        RECT 57.950 167.990 61.935 168.130 ;
        RECT 57.950 167.930 58.270 167.990 ;
        RECT 61.645 167.945 61.935 167.990 ;
        RECT 62.105 167.945 62.395 168.175 ;
        RECT 71.750 167.930 72.070 168.190 ;
        RECT 81.960 168.130 82.100 168.625 ;
        RECT 82.790 168.610 83.110 168.870 ;
        RECT 86.560 168.855 86.700 169.010 ;
        RECT 86.930 168.965 87.360 169.195 ;
        RECT 92.925 169.150 93.215 169.195 ;
        RECT 87.940 169.010 93.215 169.150 ;
        RECT 86.930 168.950 87.250 168.965 ;
        RECT 87.940 168.870 88.080 169.010 ;
        RECT 92.925 168.965 93.215 169.010 ;
        RECT 95.670 169.150 95.990 169.210 ;
        RECT 97.525 169.150 97.815 169.195 ;
        RECT 95.670 169.010 97.815 169.150 ;
        RECT 95.670 168.950 95.990 169.010 ;
        RECT 97.525 168.965 97.815 169.010 ;
        RECT 97.970 169.150 98.290 169.210 ;
        RECT 99.825 169.150 100.115 169.195 ;
        RECT 100.270 169.150 100.590 169.210 ;
        RECT 97.970 169.010 100.590 169.150 ;
        RECT 97.970 168.950 98.290 169.010 ;
        RECT 99.825 168.965 100.115 169.010 ;
        RECT 100.270 168.950 100.590 169.010 ;
        RECT 101.190 169.150 101.510 169.210 ;
        RECT 109.100 169.150 109.240 169.350 ;
        RECT 110.865 169.305 111.155 169.350 ;
        RECT 112.230 169.290 112.550 169.550 ;
        RECT 101.190 169.010 109.240 169.150 ;
        RECT 101.190 168.950 101.510 169.010 ;
        RECT 109.470 168.950 109.790 169.210 ;
        RECT 84.190 168.810 84.480 168.855 ;
        RECT 86.030 168.810 86.320 168.855 ;
        RECT 84.190 168.670 86.320 168.810 ;
        RECT 84.190 168.625 84.480 168.670 ;
        RECT 86.030 168.625 86.320 168.670 ;
        RECT 86.485 168.625 86.775 168.855 ;
        RECT 87.850 168.610 88.170 168.870 ;
        RECT 88.375 168.810 88.665 168.855 ;
        RECT 90.215 168.810 90.505 168.855 ;
        RECT 88.375 168.670 90.505 168.810 ;
        RECT 88.375 168.625 88.665 168.670 ;
        RECT 90.215 168.625 90.505 168.670 ;
        RECT 93.370 168.610 93.690 168.870 ;
        RECT 93.830 168.810 94.150 168.870 ;
        RECT 101.650 168.855 101.970 168.870 ;
        RECT 94.305 168.810 94.595 168.855 ;
        RECT 93.830 168.670 94.595 168.810 ;
        RECT 93.830 168.610 94.150 168.670 ;
        RECT 94.305 168.625 94.595 168.670 ;
        RECT 96.605 168.625 96.895 168.855 ;
        RECT 98.910 168.810 99.200 168.855 ;
        RECT 100.750 168.810 101.040 168.855 ;
        RECT 98.910 168.670 101.040 168.810 ;
        RECT 98.910 168.625 99.200 168.670 ;
        RECT 100.750 168.625 101.040 168.670 ;
        RECT 101.650 168.625 102.080 168.855 ;
        RECT 83.270 168.470 83.560 168.515 ;
        RECT 88.790 168.470 89.080 168.515 ;
        RECT 89.710 168.470 90.000 168.515 ;
        RECT 83.270 168.330 90.000 168.470 ;
        RECT 83.270 168.285 83.560 168.330 ;
        RECT 88.790 168.285 89.080 168.330 ;
        RECT 89.710 168.285 90.000 168.330 ;
        RECT 90.150 168.130 90.470 168.190 ;
        RECT 92.910 168.130 93.230 168.190 ;
        RECT 81.960 167.990 93.230 168.130 ;
        RECT 96.680 168.130 96.820 168.625 ;
        RECT 101.650 168.610 101.970 168.625 ;
        RECT 102.570 168.610 102.890 168.870 ;
        RECT 103.095 168.810 103.385 168.855 ;
        RECT 104.935 168.810 105.225 168.855 ;
        RECT 109.025 168.810 109.315 168.855 ;
        RECT 103.095 168.670 105.225 168.810 ;
        RECT 103.095 168.625 103.385 168.670 ;
        RECT 104.935 168.625 105.225 168.670 ;
        RECT 105.420 168.670 109.315 168.810 ;
        RECT 97.990 168.470 98.280 168.515 ;
        RECT 103.510 168.470 103.800 168.515 ;
        RECT 104.430 168.470 104.720 168.515 ;
        RECT 97.990 168.330 104.720 168.470 ;
        RECT 97.990 168.285 98.280 168.330 ;
        RECT 103.510 168.285 103.800 168.330 ;
        RECT 104.430 168.285 104.720 168.330 ;
        RECT 100.270 168.130 100.590 168.190 ;
        RECT 96.680 167.990 100.590 168.130 ;
        RECT 90.150 167.930 90.470 167.990 ;
        RECT 92.910 167.930 93.230 167.990 ;
        RECT 100.270 167.930 100.590 167.990 ;
        RECT 102.570 168.130 102.890 168.190 ;
        RECT 105.420 168.130 105.560 168.670 ;
        RECT 109.025 168.625 109.315 168.670 ;
        RECT 102.570 167.990 105.560 168.130 ;
        RECT 108.090 168.130 108.410 168.190 ;
        RECT 108.565 168.130 108.855 168.175 ;
        RECT 109.930 168.130 110.250 168.190 ;
        RECT 108.090 167.990 110.250 168.130 ;
        RECT 102.570 167.930 102.890 167.990 ;
        RECT 108.090 167.930 108.410 167.990 ;
        RECT 108.565 167.945 108.855 167.990 ;
        RECT 109.930 167.930 110.250 167.990 ;
        RECT 50.605 167.110 50.895 167.155 ;
        RECT 54.270 167.110 54.590 167.170 ;
        RECT 50.605 166.970 54.590 167.110 ;
        RECT 50.605 166.925 50.895 166.970 ;
        RECT 54.270 166.910 54.590 166.970 ;
        RECT 54.730 167.110 55.050 167.170 ;
        RECT 68.530 167.110 68.850 167.170 ;
        RECT 71.305 167.110 71.595 167.155 ;
        RECT 93.370 167.110 93.690 167.170 ;
        RECT 97.065 167.110 97.355 167.155 ;
        RECT 102.570 167.110 102.890 167.170 ;
        RECT 54.730 166.970 62.780 167.110 ;
        RECT 54.730 166.910 55.050 166.970 ;
        RECT 51.980 166.770 52.270 166.815 ;
        RECT 52.900 166.770 53.190 166.815 ;
        RECT 58.420 166.770 58.710 166.815 ;
        RECT 51.980 166.630 58.710 166.770 ;
        RECT 51.980 166.585 52.270 166.630 ;
        RECT 52.900 166.585 53.190 166.630 ;
        RECT 58.420 166.585 58.710 166.630 ;
        RECT 54.730 166.475 55.050 166.490 ;
        RECT 51.475 166.430 51.765 166.475 ;
        RECT 53.315 166.430 53.605 166.475 ;
        RECT 51.475 166.290 53.605 166.430 ;
        RECT 51.475 166.245 51.765 166.290 ;
        RECT 53.315 166.245 53.605 166.290 ;
        RECT 54.620 166.245 55.050 166.475 ;
        RECT 54.730 166.230 55.050 166.245 ;
        RECT 55.190 166.230 55.510 166.490 ;
        RECT 55.660 166.430 55.950 166.475 ;
        RECT 57.500 166.430 57.790 166.475 ;
        RECT 59.115 166.430 59.405 166.475 ;
        RECT 55.660 166.290 57.790 166.430 ;
        RECT 55.660 166.245 55.950 166.290 ;
        RECT 57.500 166.245 57.790 166.290 ;
        RECT 58.500 166.290 59.405 166.430 ;
        RECT 62.640 166.430 62.780 166.970 ;
        RECT 68.530 166.970 71.595 167.110 ;
        RECT 68.530 166.910 68.850 166.970 ;
        RECT 71.305 166.925 71.595 166.970 ;
        RECT 72.300 166.970 79.800 167.110 ;
        RECT 71.750 166.570 72.070 166.830 ;
        RECT 72.300 166.430 72.440 166.970 ;
        RECT 76.825 166.770 77.115 166.815 ;
        RECT 77.730 166.770 78.050 166.830 ;
        RECT 76.825 166.630 78.050 166.770 ;
        RECT 76.825 166.585 77.115 166.630 ;
        RECT 77.730 166.570 78.050 166.630 ;
        RECT 62.640 166.290 72.440 166.430 ;
        RECT 75.430 166.430 75.750 166.490 ;
        RECT 79.660 166.475 79.800 166.970 ;
        RECT 93.370 166.970 102.890 167.110 ;
        RECT 93.370 166.910 93.690 166.970 ;
        RECT 97.065 166.925 97.355 166.970 ;
        RECT 102.570 166.910 102.890 166.970 ;
        RECT 103.950 166.910 104.270 167.170 ;
        RECT 104.885 167.110 105.175 167.155 ;
        RECT 109.470 167.110 109.790 167.170 ;
        RECT 104.885 166.970 109.790 167.110 ;
        RECT 104.885 166.925 105.175 166.970 ;
        RECT 109.470 166.910 109.790 166.970 ;
        RECT 80.490 166.570 80.810 166.830 ;
        RECT 104.040 166.770 104.180 166.910 ;
        RECT 111.770 166.770 112.090 166.830 ;
        RECT 92.080 166.630 95.900 166.770 ;
        RECT 104.040 166.630 112.090 166.770 ;
        RECT 92.080 166.490 92.220 166.630 ;
        RECT 75.905 166.430 76.195 166.475 ;
        RECT 75.430 166.290 76.195 166.430 ;
        RECT 58.500 166.150 58.640 166.290 ;
        RECT 59.115 166.245 59.405 166.290 ;
        RECT 75.430 166.230 75.750 166.290 ;
        RECT 75.905 166.245 76.195 166.290 ;
        RECT 79.585 166.430 79.875 166.475 ;
        RECT 81.410 166.430 81.730 166.490 ;
        RECT 79.585 166.290 81.730 166.430 ;
        RECT 79.585 166.245 79.875 166.290 ;
        RECT 81.410 166.230 81.730 166.290 ;
        RECT 91.990 166.230 92.310 166.490 ;
        RECT 92.450 166.230 92.770 166.490 ;
        RECT 93.830 166.230 94.150 166.490 ;
        RECT 95.760 166.475 95.900 166.630 ;
        RECT 111.770 166.570 112.090 166.630 ;
        RECT 94.765 166.245 95.055 166.475 ;
        RECT 95.685 166.245 95.975 166.475 ;
        RECT 96.130 166.430 96.450 166.490 ;
        RECT 101.650 166.430 101.970 166.490 ;
        RECT 96.130 166.290 101.970 166.430 ;
        RECT 53.810 165.890 54.130 166.150 ;
        RECT 58.410 165.890 58.730 166.150 ;
        RECT 59.790 165.890 60.110 166.150 ;
        RECT 77.745 166.090 78.035 166.135 ;
        RECT 93.920 166.090 94.060 166.230 ;
        RECT 77.745 165.950 94.060 166.090 ;
        RECT 77.745 165.905 78.035 165.950 ;
        RECT 94.305 165.905 94.595 166.135 ;
        RECT 52.395 165.750 52.685 165.795 ;
        RECT 55.625 165.750 55.915 165.795 ;
        RECT 52.395 165.610 55.915 165.750 ;
        RECT 52.395 165.565 52.685 165.610 ;
        RECT 55.625 165.565 55.915 165.610 ;
        RECT 56.585 165.750 56.875 165.795 ;
        RECT 57.490 165.750 57.810 165.810 ;
        RECT 74.985 165.750 75.275 165.795 ;
        RECT 91.545 165.750 91.835 165.795 ;
        RECT 94.380 165.750 94.520 165.905 ;
        RECT 56.585 165.610 57.810 165.750 ;
        RECT 56.585 165.565 56.875 165.610 ;
        RECT 57.490 165.550 57.810 165.610 ;
        RECT 61.260 165.610 94.520 165.750 ;
        RECT 59.790 165.410 60.110 165.470 ;
        RECT 61.260 165.410 61.400 165.610 ;
        RECT 74.985 165.565 75.275 165.610 ;
        RECT 91.545 165.565 91.835 165.610 ;
        RECT 59.790 165.270 61.400 165.410 ;
        RECT 72.670 165.410 72.990 165.470 ;
        RECT 94.840 165.410 94.980 166.245 ;
        RECT 96.130 166.230 96.450 166.290 ;
        RECT 101.650 166.230 101.970 166.290 ;
        RECT 103.950 166.430 104.270 166.490 ;
        RECT 105.330 166.430 105.650 166.490 ;
        RECT 107.185 166.430 107.475 166.475 ;
        RECT 110.850 166.430 111.170 166.490 ;
        RECT 112.245 166.430 112.535 166.475 ;
        RECT 103.950 166.290 105.100 166.430 ;
        RECT 103.950 166.230 104.270 166.290 ;
        RECT 104.410 165.890 104.730 166.150 ;
        RECT 104.960 166.090 105.100 166.290 ;
        RECT 105.330 166.290 107.475 166.430 ;
        RECT 105.330 166.230 105.650 166.290 ;
        RECT 107.185 166.245 107.475 166.290 ;
        RECT 107.720 166.290 112.535 166.430 ;
        RECT 107.720 166.090 107.860 166.290 ;
        RECT 110.850 166.230 111.170 166.290 ;
        RECT 112.245 166.245 112.535 166.290 ;
        RECT 104.960 165.950 107.860 166.090 ;
        RECT 108.090 165.890 108.410 166.150 ;
        RECT 112.705 165.905 112.995 166.135 ;
        RECT 103.490 165.550 103.810 165.810 ;
        RECT 104.500 165.750 104.640 165.890 ;
        RECT 111.310 165.750 111.630 165.810 ;
        RECT 112.780 165.750 112.920 165.905 ;
        RECT 104.500 165.610 112.920 165.750 ;
        RECT 111.310 165.550 111.630 165.610 ;
        RECT 96.590 165.410 96.910 165.470 ;
        RECT 72.670 165.270 96.910 165.410 ;
        RECT 103.580 165.410 103.720 165.550 ;
        RECT 106.725 165.410 107.015 165.455 ;
        RECT 103.580 165.270 107.015 165.410 ;
        RECT 59.790 165.210 60.110 165.270 ;
        RECT 72.670 165.210 72.990 165.270 ;
        RECT 96.590 165.210 96.910 165.270 ;
        RECT 106.725 165.225 107.015 165.270 ;
        RECT 109.930 165.210 110.250 165.470 ;
        RECT 61.185 164.390 61.475 164.435 ;
        RECT 63.470 164.390 63.790 164.450 ;
        RECT 82.330 164.390 82.650 164.450 ;
        RECT 61.185 164.250 63.790 164.390 ;
        RECT 61.185 164.205 61.475 164.250 ;
        RECT 63.470 164.190 63.790 164.250 ;
        RECT 66.780 164.250 82.650 164.390 ;
        RECT 62.975 164.050 63.265 164.095 ;
        RECT 66.205 164.050 66.495 164.095 ;
        RECT 62.975 163.910 66.495 164.050 ;
        RECT 62.975 163.865 63.265 163.910 ;
        RECT 66.205 163.865 66.495 163.910 ;
        RECT 55.190 163.710 55.510 163.770 ;
        RECT 56.585 163.710 56.875 163.755 ;
        RECT 64.405 163.710 64.695 163.755 ;
        RECT 66.780 163.710 66.920 164.250 ;
        RECT 82.330 164.190 82.650 164.250 ;
        RECT 84.185 164.390 84.475 164.435 ;
        RECT 86.470 164.390 86.790 164.450 ;
        RECT 84.185 164.250 86.790 164.390 ;
        RECT 84.185 164.205 84.475 164.250 ;
        RECT 86.470 164.190 86.790 164.250 ;
        RECT 92.450 164.390 92.770 164.450 ;
        RECT 93.845 164.390 94.135 164.435 ;
        RECT 92.450 164.250 94.135 164.390 ;
        RECT 92.450 164.190 92.770 164.250 ;
        RECT 93.845 164.205 94.135 164.250 ;
        RECT 96.590 164.390 96.910 164.450 ;
        RECT 103.030 164.390 103.350 164.450 ;
        RECT 96.590 164.250 103.350 164.390 ;
        RECT 96.590 164.190 96.910 164.250 ;
        RECT 103.030 164.190 103.350 164.250 ;
        RECT 112.245 164.390 112.535 164.435 ;
        RECT 116.830 164.390 117.150 164.450 ;
        RECT 112.245 164.250 117.150 164.390 ;
        RECT 112.245 164.205 112.535 164.250 ;
        RECT 116.830 164.190 117.150 164.250 ;
        RECT 67.150 163.850 67.470 164.110 ;
        RECT 70.830 164.050 71.150 164.110 ;
        RECT 68.160 163.910 71.150 164.050 ;
        RECT 55.190 163.570 56.875 163.710 ;
        RECT 55.190 163.510 55.510 163.570 ;
        RECT 56.585 163.525 56.875 163.570 ;
        RECT 60.800 163.570 66.920 163.710 ;
        RECT 67.240 163.710 67.380 163.850 ;
        RECT 68.160 163.710 68.300 163.910 ;
        RECT 70.830 163.850 71.150 163.910 ;
        RECT 74.970 164.050 75.290 164.110 ;
        RECT 82.790 164.050 83.110 164.110 ;
        RECT 104.410 164.050 104.730 164.110 ;
        RECT 74.970 163.910 88.080 164.050 ;
        RECT 74.970 163.850 75.290 163.910 ;
        RECT 82.790 163.850 83.110 163.910 ;
        RECT 67.240 163.570 68.300 163.710 ;
        RECT 69.450 163.710 69.770 163.770 ;
        RECT 73.130 163.710 73.450 163.770 ;
        RECT 69.450 163.570 73.450 163.710 ;
        RECT 57.045 163.370 57.335 163.415 ;
        RECT 59.790 163.370 60.110 163.430 ;
        RECT 57.045 163.230 60.110 163.370 ;
        RECT 57.045 163.185 57.335 163.230 ;
        RECT 59.790 163.170 60.110 163.230 ;
        RECT 53.810 163.030 54.130 163.090 ;
        RECT 60.800 163.030 60.940 163.570 ;
        RECT 64.405 163.525 64.695 163.570 ;
        RECT 69.450 163.510 69.770 163.570 ;
        RECT 73.130 163.510 73.450 163.570 ;
        RECT 79.200 163.570 82.100 163.710 ;
        RECT 65.310 163.415 65.630 163.430 ;
        RECT 62.055 163.370 62.345 163.415 ;
        RECT 63.895 163.370 64.185 163.415 ;
        RECT 62.055 163.230 64.185 163.370 ;
        RECT 62.055 163.185 62.345 163.230 ;
        RECT 63.895 163.185 64.185 163.230 ;
        RECT 65.200 163.185 65.630 163.415 ;
        RECT 65.310 163.170 65.630 163.185 ;
        RECT 65.770 163.170 66.090 163.430 ;
        RECT 66.240 163.370 66.530 163.415 ;
        RECT 68.080 163.370 68.370 163.415 ;
        RECT 66.240 163.230 68.370 163.370 ;
        RECT 66.240 163.185 66.530 163.230 ;
        RECT 68.080 163.185 68.370 163.230 ;
        RECT 69.910 163.370 70.230 163.430 ;
        RECT 70.385 163.370 70.675 163.415 ;
        RECT 72.670 163.370 72.990 163.430 ;
        RECT 69.910 163.230 72.990 163.370 ;
        RECT 69.910 163.170 70.230 163.230 ;
        RECT 70.385 163.185 70.675 163.230 ;
        RECT 72.670 163.170 72.990 163.230 ;
        RECT 53.810 162.890 60.940 163.030 ;
        RECT 62.560 163.030 62.850 163.075 ;
        RECT 63.480 163.030 63.770 163.075 ;
        RECT 69.000 163.030 69.290 163.075 ;
        RECT 62.560 162.890 69.290 163.030 ;
        RECT 53.810 162.830 54.130 162.890 ;
        RECT 62.560 162.845 62.850 162.890 ;
        RECT 63.480 162.845 63.770 162.890 ;
        RECT 69.000 162.845 69.290 162.890 ;
        RECT 55.190 162.490 55.510 162.750 ;
        RECT 65.310 162.690 65.630 162.750 ;
        RECT 77.730 162.690 78.050 162.750 ;
        RECT 79.200 162.735 79.340 163.570 ;
        RECT 81.410 163.170 81.730 163.430 ;
        RECT 81.960 163.415 82.100 163.570 ;
        RECT 81.885 163.185 82.175 163.415 ;
        RECT 82.330 163.370 82.650 163.430 ;
        RECT 82.805 163.370 83.095 163.415 ;
        RECT 85.090 163.370 85.410 163.430 ;
        RECT 87.940 163.415 88.080 163.910 ;
        RECT 100.820 163.910 104.730 164.050 ;
        RECT 88.785 163.710 89.075 163.755 ;
        RECT 89.690 163.710 90.010 163.770 ;
        RECT 88.785 163.570 90.010 163.710 ;
        RECT 88.785 163.525 89.075 163.570 ;
        RECT 89.690 163.510 90.010 163.570 ;
        RECT 90.150 163.510 90.470 163.770 ;
        RECT 94.750 163.710 95.070 163.770 ;
        RECT 100.820 163.755 100.960 163.910 ;
        RECT 104.410 163.850 104.730 163.910 ;
        RECT 105.790 164.050 106.110 164.110 ;
        RECT 107.170 164.050 107.490 164.110 ;
        RECT 109.485 164.050 109.775 164.095 ;
        RECT 105.790 163.910 109.775 164.050 ;
        RECT 105.790 163.850 106.110 163.910 ;
        RECT 107.170 163.850 107.490 163.910 ;
        RECT 109.485 163.865 109.775 163.910 ;
        RECT 96.605 163.710 96.895 163.755 ;
        RECT 100.745 163.710 101.035 163.755 ;
        RECT 94.750 163.570 101.035 163.710 ;
        RECT 94.750 163.510 95.070 163.570 ;
        RECT 96.605 163.525 96.895 163.570 ;
        RECT 100.745 163.525 101.035 163.570 ;
        RECT 101.190 163.510 101.510 163.770 ;
        RECT 82.330 163.230 85.410 163.370 ;
        RECT 82.330 163.170 82.650 163.230 ;
        RECT 82.805 163.185 83.095 163.230 ;
        RECT 85.090 163.170 85.410 163.230 ;
        RECT 87.865 163.185 88.155 163.415 ;
        RECT 88.325 163.370 88.615 163.415 ;
        RECT 90.240 163.370 90.380 163.510 ;
        RECT 88.325 163.230 90.380 163.370 ;
        RECT 88.325 163.185 88.615 163.230 ;
        RECT 95.210 163.170 95.530 163.430 ;
        RECT 96.145 163.370 96.435 163.415 ;
        RECT 101.280 163.370 101.420 163.510 ;
        RECT 96.145 163.230 101.420 163.370 ;
        RECT 109.930 163.370 110.250 163.430 ;
        RECT 110.405 163.370 110.695 163.415 ;
        RECT 109.930 163.230 110.695 163.370 ;
        RECT 96.145 163.185 96.435 163.230 ;
        RECT 109.930 163.170 110.250 163.230 ;
        RECT 110.405 163.185 110.695 163.230 ;
        RECT 79.585 163.030 79.875 163.075 ;
        RECT 79.585 162.890 86.240 163.030 ;
        RECT 79.585 162.845 79.875 162.890 ;
        RECT 86.100 162.735 86.240 162.890 ;
        RECT 89.230 162.830 89.550 163.090 ;
        RECT 95.300 163.030 95.440 163.170 ;
        RECT 99.825 163.030 100.115 163.075 ;
        RECT 101.190 163.030 101.510 163.090 ;
        RECT 95.300 162.890 101.510 163.030 ;
        RECT 99.825 162.845 100.115 162.890 ;
        RECT 101.190 162.830 101.510 162.890 ;
        RECT 102.570 162.830 102.890 163.090 ;
        RECT 103.950 163.030 104.270 163.090 ;
        RECT 103.950 162.890 111.080 163.030 ;
        RECT 103.950 162.830 104.270 162.890 ;
        RECT 79.125 162.690 79.415 162.735 ;
        RECT 65.310 162.550 79.415 162.690 ;
        RECT 65.310 162.490 65.630 162.550 ;
        RECT 77.730 162.490 78.050 162.550 ;
        RECT 79.125 162.505 79.415 162.550 ;
        RECT 86.025 162.505 86.315 162.735 ;
        RECT 89.320 162.690 89.460 162.830 ;
        RECT 95.685 162.690 95.975 162.735 ;
        RECT 96.130 162.690 96.450 162.750 ;
        RECT 89.320 162.550 96.450 162.690 ;
        RECT 95.685 162.505 95.975 162.550 ;
        RECT 96.130 162.490 96.450 162.550 ;
        RECT 97.985 162.690 98.275 162.735 ;
        RECT 98.430 162.690 98.750 162.750 ;
        RECT 97.985 162.550 98.750 162.690 ;
        RECT 97.985 162.505 98.275 162.550 ;
        RECT 98.430 162.490 98.750 162.550 ;
        RECT 99.350 162.690 99.670 162.750 ;
        RECT 100.285 162.690 100.575 162.735 ;
        RECT 109.010 162.690 109.330 162.750 ;
        RECT 110.940 162.735 111.080 162.890 ;
        RECT 99.350 162.550 109.330 162.690 ;
        RECT 99.350 162.490 99.670 162.550 ;
        RECT 100.285 162.505 100.575 162.550 ;
        RECT 109.010 162.490 109.330 162.550 ;
        RECT 110.865 162.505 111.155 162.735 ;
        RECT 54.730 161.470 55.050 161.730 ;
        RECT 57.950 161.470 58.270 161.730 ;
        RECT 65.310 161.670 65.630 161.730 ;
        RECT 62.180 161.530 65.630 161.670 ;
        RECT 54.820 161.330 54.960 161.470 ;
        RECT 53.440 161.190 54.960 161.330 ;
        RECT 52.890 160.790 53.210 161.050 ;
        RECT 53.440 160.695 53.580 161.190 ;
        RECT 62.180 161.035 62.320 161.530 ;
        RECT 65.310 161.470 65.630 161.530 ;
        RECT 69.925 161.670 70.215 161.715 ;
        RECT 70.370 161.670 70.690 161.730 ;
        RECT 69.925 161.530 70.690 161.670 ;
        RECT 69.925 161.485 70.215 161.530 ;
        RECT 70.370 161.470 70.690 161.530 ;
        RECT 73.590 161.670 73.910 161.730 ;
        RECT 74.065 161.670 74.355 161.715 ;
        RECT 73.590 161.530 74.355 161.670 ;
        RECT 73.590 161.470 73.910 161.530 ;
        RECT 74.065 161.485 74.355 161.530 ;
        RECT 75.905 161.670 76.195 161.715 ;
        RECT 76.350 161.670 76.670 161.730 ;
        RECT 75.905 161.530 76.670 161.670 ;
        RECT 75.905 161.485 76.195 161.530 ;
        RECT 76.350 161.470 76.670 161.530 ;
        RECT 98.430 161.470 98.750 161.730 ;
        RECT 101.665 161.670 101.955 161.715 ;
        RECT 102.570 161.670 102.890 161.730 ;
        RECT 101.665 161.530 102.890 161.670 ;
        RECT 101.665 161.485 101.955 161.530 ;
        RECT 102.570 161.470 102.890 161.530 ;
        RECT 103.030 161.670 103.350 161.730 ;
        RECT 105.330 161.670 105.650 161.730 ;
        RECT 105.805 161.670 106.095 161.715 ;
        RECT 103.030 161.530 104.640 161.670 ;
        RECT 103.030 161.470 103.350 161.530 ;
        RECT 65.770 161.330 66.090 161.390 ;
        RECT 62.640 161.190 66.090 161.330 ;
        RECT 56.125 160.990 56.415 161.035 ;
        RECT 54.820 160.850 56.415 160.990 ;
        RECT 54.820 160.695 54.960 160.850 ;
        RECT 56.125 160.805 56.415 160.850 ;
        RECT 62.105 160.805 62.395 161.035 ;
        RECT 53.365 160.465 53.655 160.695 ;
        RECT 54.745 160.465 55.035 160.695 ;
        RECT 55.190 160.650 55.510 160.710 ;
        RECT 62.640 160.695 62.780 161.190 ;
        RECT 65.770 161.130 66.090 161.190 ;
        RECT 76.810 161.330 77.130 161.390 ;
        RECT 96.605 161.330 96.895 161.375 ;
        RECT 98.520 161.330 98.660 161.470 ;
        RECT 76.810 161.190 79.800 161.330 ;
        RECT 76.810 161.130 77.130 161.190 ;
        RECT 65.325 160.990 65.615 161.035 ;
        RECT 69.450 160.990 69.770 161.050 ;
        RECT 65.325 160.850 69.770 160.990 ;
        RECT 65.325 160.805 65.615 160.850 ;
        RECT 69.450 160.790 69.770 160.850 ;
        RECT 71.765 160.990 72.055 161.035 ;
        RECT 74.970 160.990 75.290 161.050 ;
        RECT 71.765 160.850 75.290 160.990 ;
        RECT 71.765 160.805 72.055 160.850 ;
        RECT 74.970 160.790 75.290 160.850 ;
        RECT 55.665 160.650 55.955 160.695 ;
        RECT 55.190 160.510 55.955 160.650 ;
        RECT 55.190 160.450 55.510 160.510 ;
        RECT 55.665 160.465 55.955 160.510 ;
        RECT 62.565 160.465 62.855 160.695 ;
        RECT 65.785 160.650 66.075 160.695 ;
        RECT 69.910 160.650 70.230 160.710 ;
        RECT 65.785 160.510 70.230 160.650 ;
        RECT 65.785 160.465 66.075 160.510 ;
        RECT 69.910 160.450 70.230 160.510 ;
        RECT 72.210 160.450 72.530 160.710 ;
        RECT 73.145 160.650 73.435 160.695 ;
        RECT 74.050 160.650 74.370 160.710 ;
        RECT 73.145 160.510 74.370 160.650 ;
        RECT 73.145 160.465 73.435 160.510 ;
        RECT 74.050 160.450 74.370 160.510 ;
        RECT 76.350 160.450 76.670 160.710 ;
        RECT 79.660 160.695 79.800 161.190 ;
        RECT 96.605 161.190 98.660 161.330 ;
        RECT 100.270 161.330 100.590 161.390 ;
        RECT 103.950 161.330 104.270 161.390 ;
        RECT 100.270 161.190 104.270 161.330 ;
        RECT 104.500 161.330 104.640 161.530 ;
        RECT 105.330 161.530 106.095 161.670 ;
        RECT 105.330 161.470 105.650 161.530 ;
        RECT 105.805 161.485 106.095 161.530 ;
        RECT 110.850 161.470 111.170 161.730 ;
        RECT 112.230 161.470 112.550 161.730 ;
        RECT 106.725 161.330 107.015 161.375 ;
        RECT 104.500 161.190 107.015 161.330 ;
        RECT 96.605 161.145 96.895 161.190 ;
        RECT 100.270 161.130 100.590 161.190 ;
        RECT 103.950 161.130 104.270 161.190 ;
        RECT 106.725 161.145 107.015 161.190 ;
        RECT 80.045 160.990 80.335 161.035 ;
        RECT 82.330 160.990 82.650 161.050 ;
        RECT 80.045 160.850 82.650 160.990 ;
        RECT 80.045 160.805 80.335 160.850 ;
        RECT 82.330 160.790 82.650 160.850 ;
        RECT 91.530 160.790 91.850 161.050 ;
        RECT 103.505 160.990 103.795 161.035 ;
        RECT 99.900 160.850 103.795 160.990 ;
        RECT 76.825 160.465 77.115 160.695 ;
        RECT 79.585 160.465 79.875 160.695 ;
        RECT 63.945 160.310 64.235 160.355 ;
        RECT 67.610 160.310 67.930 160.370 ;
        RECT 63.945 160.170 67.930 160.310 ;
        RECT 74.140 160.310 74.280 160.450 ;
        RECT 76.900 160.310 77.040 160.465 ;
        RECT 91.990 160.450 92.310 160.710 ;
        RECT 96.130 160.650 96.450 160.710 ;
        RECT 99.900 160.650 100.040 160.850 ;
        RECT 103.505 160.805 103.795 160.850 ;
        RECT 96.130 160.510 100.040 160.650 ;
        RECT 96.130 160.450 96.450 160.510 ;
        RECT 104.410 160.450 104.730 160.710 ;
        RECT 104.870 160.650 105.190 160.710 ;
        RECT 107.645 160.650 107.935 160.695 ;
        RECT 104.870 160.510 107.935 160.650 ;
        RECT 104.870 160.450 105.190 160.510 ;
        RECT 107.645 160.465 107.935 160.510 ;
        RECT 95.685 160.310 95.975 160.355 ;
        RECT 108.550 160.310 108.870 160.370 ;
        RECT 74.140 160.170 77.040 160.310 ;
        RECT 81.040 160.170 108.870 160.310 ;
        RECT 63.945 160.125 64.235 160.170 ;
        RECT 67.610 160.110 67.930 160.170 ;
        RECT 81.040 160.030 81.180 160.170 ;
        RECT 95.685 160.125 95.975 160.170 ;
        RECT 108.550 160.110 108.870 160.170 ;
        RECT 67.150 159.770 67.470 160.030 ;
        RECT 80.950 159.770 81.270 160.030 ;
        RECT 81.410 159.770 81.730 160.030 ;
        RECT 89.690 159.770 90.010 160.030 ;
        RECT 44.610 158.750 44.930 159.010 ;
        RECT 56.110 158.750 56.430 159.010 ;
        RECT 59.805 158.950 60.095 158.995 ;
        RECT 61.630 158.950 61.950 159.010 ;
        RECT 59.805 158.810 61.950 158.950 ;
        RECT 59.805 158.765 60.095 158.810 ;
        RECT 61.630 158.750 61.950 158.810 ;
        RECT 64.390 158.950 64.710 159.010 ;
        RECT 64.865 158.950 65.155 158.995 ;
        RECT 64.390 158.810 65.155 158.950 ;
        RECT 64.390 158.750 64.710 158.810 ;
        RECT 64.865 158.765 65.155 158.810 ;
        RECT 67.150 158.750 67.470 159.010 ;
        RECT 67.610 158.750 67.930 159.010 ;
        RECT 70.385 158.950 70.675 158.995 ;
        RECT 72.210 158.950 72.530 159.010 ;
        RECT 70.385 158.810 72.530 158.950 ;
        RECT 70.385 158.765 70.675 158.810 ;
        RECT 72.210 158.750 72.530 158.810 ;
        RECT 74.970 158.750 75.290 159.010 ;
        RECT 77.270 158.950 77.590 159.010 ;
        RECT 79.125 158.950 79.415 158.995 ;
        RECT 77.270 158.810 79.415 158.950 ;
        RECT 77.270 158.750 77.590 158.810 ;
        RECT 79.125 158.765 79.415 158.810 ;
        RECT 81.410 158.750 81.730 159.010 ;
        RECT 87.405 158.950 87.695 158.995 ;
        RECT 89.230 158.950 89.550 159.010 ;
        RECT 87.405 158.810 89.550 158.950 ;
        RECT 87.405 158.765 87.695 158.810 ;
        RECT 89.230 158.750 89.550 158.810 ;
        RECT 89.690 158.750 90.010 159.010 ;
        RECT 90.165 158.950 90.455 158.995 ;
        RECT 90.610 158.950 90.930 159.010 ;
        RECT 90.165 158.810 90.930 158.950 ;
        RECT 90.165 158.765 90.455 158.810 ;
        RECT 90.610 158.750 90.930 158.810 ;
        RECT 95.225 158.950 95.515 158.995 ;
        RECT 95.670 158.950 95.990 159.010 ;
        RECT 95.225 158.810 95.990 158.950 ;
        RECT 95.225 158.765 95.515 158.810 ;
        RECT 95.670 158.750 95.990 158.810 ;
        RECT 100.285 158.950 100.575 158.995 ;
        RECT 100.730 158.950 101.050 159.010 ;
        RECT 100.285 158.810 101.050 158.950 ;
        RECT 100.285 158.765 100.575 158.810 ;
        RECT 100.730 158.750 101.050 158.810 ;
        RECT 101.190 158.950 101.510 159.010 ;
        RECT 105.345 158.950 105.635 158.995 ;
        RECT 101.190 158.810 105.635 158.950 ;
        RECT 101.190 158.750 101.510 158.810 ;
        RECT 105.345 158.765 105.635 158.810 ;
        RECT 108.090 158.950 108.410 159.010 ;
        RECT 109.945 158.950 110.235 158.995 ;
        RECT 108.090 158.810 110.235 158.950 ;
        RECT 108.090 158.750 108.410 158.810 ;
        RECT 109.945 158.765 110.235 158.810 ;
        RECT 111.770 158.950 112.090 159.010 ;
        RECT 113.165 158.950 113.455 158.995 ;
        RECT 111.770 158.810 113.455 158.950 ;
        RECT 111.770 158.750 112.090 158.810 ;
        RECT 113.165 158.765 113.455 158.810 ;
        RECT 49.685 158.610 49.975 158.655 ;
        RECT 62.550 158.610 62.870 158.670 ;
        RECT 49.685 158.470 62.870 158.610 ;
        RECT 49.685 158.425 49.975 158.470 ;
        RECT 62.550 158.410 62.870 158.470 ;
        RECT 52.890 158.070 53.210 158.330 ;
        RECT 43.690 157.730 44.010 157.990 ;
        RECT 48.750 157.730 49.070 157.990 ;
        RECT 52.980 157.590 53.120 158.070 ;
        RECT 53.350 157.930 53.670 157.990 ;
        RECT 55.205 157.930 55.495 157.975 ;
        RECT 53.350 157.790 55.495 157.930 ;
        RECT 53.350 157.730 53.670 157.790 ;
        RECT 55.205 157.745 55.495 157.790 ;
        RECT 58.870 157.730 59.190 157.990 ;
        RECT 63.930 157.730 64.250 157.990 ;
        RECT 67.240 157.930 67.380 158.750 ;
        RECT 67.700 158.270 67.840 158.750 ;
        RECT 68.545 158.270 68.835 158.315 ;
        RECT 80.950 158.270 81.270 158.330 ;
        RECT 67.700 158.130 68.835 158.270 ;
        RECT 68.545 158.085 68.835 158.130 ;
        RECT 71.840 158.130 81.270 158.270 ;
        RECT 81.500 158.270 81.640 158.750 ;
        RECT 84.645 158.270 84.935 158.315 ;
        RECT 89.780 158.270 89.920 158.750 ;
        RECT 108.550 158.410 108.870 158.670 ;
        RECT 81.500 158.130 84.935 158.270 ;
        RECT 69.005 157.930 69.295 157.975 ;
        RECT 67.240 157.790 69.295 157.930 ;
        RECT 69.005 157.745 69.295 157.790 ;
        RECT 69.910 157.930 70.230 157.990 ;
        RECT 71.305 157.930 71.595 157.975 ;
        RECT 69.910 157.790 71.595 157.930 ;
        RECT 69.910 157.730 70.230 157.790 ;
        RECT 71.305 157.745 71.595 157.790 ;
        RECT 71.840 157.590 71.980 158.130 ;
        RECT 80.950 158.070 81.270 158.130 ;
        RECT 84.645 158.085 84.935 158.130 ;
        RECT 85.180 158.130 89.920 158.270 ;
        RECT 108.640 158.270 108.780 158.410 ;
        RECT 109.485 158.270 109.775 158.315 ;
        RECT 108.640 158.130 109.775 158.270 ;
        RECT 74.050 157.730 74.370 157.990 ;
        RECT 75.890 157.730 76.210 157.990 ;
        RECT 76.350 157.730 76.670 157.990 ;
        RECT 80.030 157.730 80.350 157.990 ;
        RECT 85.180 157.975 85.320 158.130 ;
        RECT 109.485 158.085 109.775 158.130 ;
        RECT 85.105 157.745 85.395 157.975 ;
        RECT 86.485 157.745 86.775 157.975 ;
        RECT 75.980 157.590 76.120 157.730 ;
        RECT 52.980 157.450 71.980 157.590 ;
        RECT 72.300 157.450 76.120 157.590 ;
        RECT 72.300 157.295 72.440 157.450 ;
        RECT 72.225 157.065 72.515 157.295 ;
        RECT 76.440 157.250 76.580 157.730 ;
        RECT 83.710 157.590 84.030 157.650 ;
        RECT 86.560 157.590 86.700 157.745 ;
        RECT 89.230 157.730 89.550 157.990 ;
        RECT 91.530 157.730 91.850 157.990 ;
        RECT 94.290 157.730 94.610 157.990 ;
        RECT 99.350 157.730 99.670 157.990 ;
        RECT 104.410 157.730 104.730 157.990 ;
        RECT 107.630 157.730 107.950 157.990 ;
        RECT 108.565 157.745 108.855 157.975 ;
        RECT 109.010 157.930 109.330 157.990 ;
        RECT 110.865 157.930 111.155 157.975 ;
        RECT 109.010 157.790 111.155 157.930 ;
        RECT 83.710 157.450 86.700 157.590 ;
        RECT 91.620 157.590 91.760 157.730 ;
        RECT 108.640 157.590 108.780 157.745 ;
        RECT 109.010 157.730 109.330 157.790 ;
        RECT 110.865 157.745 111.155 157.790 ;
        RECT 114.070 157.730 114.390 157.990 ;
        RECT 113.610 157.590 113.930 157.650 ;
        RECT 91.620 157.450 113.930 157.590 ;
        RECT 83.710 157.390 84.030 157.450 ;
        RECT 113.610 157.390 113.930 157.450 ;
        RECT 83.265 157.250 83.555 157.295 ;
        RECT 76.440 157.110 83.555 157.250 ;
        RECT 83.265 157.065 83.555 157.110 ;
        RECT 111.785 157.250 112.075 157.295 ;
        RECT 114.530 157.250 114.850 157.310 ;
        RECT 111.785 157.110 114.850 157.250 ;
        RECT 111.785 157.065 112.075 157.110 ;
        RECT 114.530 157.050 114.850 157.110 ;
        RECT 79.110 156.230 79.430 156.290 ;
        RECT 80.030 156.230 80.350 156.290 ;
        RECT 79.110 156.090 80.350 156.230 ;
        RECT 79.110 156.030 79.430 156.090 ;
        RECT 80.030 156.030 80.350 156.090 ;
        RECT 78.910 128.595 79.230 128.600 ;
        RECT 101.555 128.595 101.875 128.600 ;
        RECT 78.910 128.345 101.875 128.595 ;
        RECT 78.910 128.340 79.230 128.345 ;
        RECT 101.555 128.340 101.875 128.345 ;
        RECT 62.930 127.920 63.830 127.970 ;
        RECT 64.810 127.920 65.710 127.970 ;
        RECT 62.900 127.690 63.860 127.920 ;
        RECT 64.780 127.895 65.740 127.920 ;
        RECT 64.780 127.690 66.000 127.895 ;
        RECT 66.660 127.690 67.620 127.920 ;
        RECT 68.540 127.690 69.500 127.920 ;
        RECT 70.400 127.690 71.400 128.010 ;
        RECT 72.280 127.690 73.280 128.010 ;
        RECT 74.160 127.920 75.160 128.010 ;
        RECT 85.590 127.920 86.490 127.970 ;
        RECT 87.470 127.920 88.370 127.970 ;
        RECT 74.160 127.690 75.420 127.920 ;
        RECT 85.560 127.690 86.520 127.920 ;
        RECT 87.440 127.895 88.400 127.920 ;
        RECT 87.440 127.690 88.660 127.895 ;
        RECT 89.320 127.690 90.280 127.920 ;
        RECT 91.200 127.690 92.160 127.920 ;
        RECT 93.060 127.690 94.060 128.010 ;
        RECT 94.940 127.690 95.940 128.010 ;
        RECT 96.820 127.920 97.820 128.010 ;
        RECT 108.250 127.920 109.150 127.970 ;
        RECT 110.130 127.920 111.030 127.970 ;
        RECT 96.820 127.690 98.080 127.920 ;
        RECT 108.220 127.690 109.180 127.920 ;
        RECT 110.100 127.895 111.060 127.920 ;
        RECT 110.100 127.690 111.320 127.895 ;
        RECT 111.980 127.690 112.940 127.920 ;
        RECT 113.860 127.690 114.820 127.920 ;
        RECT 115.720 127.690 116.720 128.010 ;
        RECT 117.600 127.690 118.600 128.010 ;
        RECT 119.480 127.920 120.480 128.010 ;
        RECT 119.480 127.690 120.740 127.920 ;
        RECT 62.930 127.650 63.830 127.690 ;
        RECT 64.810 127.650 66.000 127.690 ;
        RECT 62.620 125.765 62.850 127.530 ;
        RECT 62.535 125.530 62.850 125.765 ;
        RECT 62.535 124.440 62.725 125.530 ;
        RECT 63.285 125.370 63.475 127.650 ;
        RECT 65.160 127.530 66.000 127.650 ;
        RECT 65.160 127.300 66.020 127.530 ;
        RECT 65.165 125.770 65.355 127.300 ;
        RECT 65.790 125.775 66.020 127.300 ;
        RECT 66.380 125.785 66.610 127.530 ;
        RECT 65.790 125.770 66.115 125.775 ;
        RECT 65.165 125.370 66.115 125.770 ;
        RECT 62.900 124.600 63.860 125.370 ;
        RECT 58.860 123.815 59.190 124.220 ;
        RECT 59.460 123.815 59.790 124.220 ;
        RECT 60.060 123.815 60.390 124.220 ;
        RECT 60.660 123.815 60.990 124.220 ;
        RECT 62.535 124.200 62.850 124.440 ;
        RECT 57.535 123.565 60.990 123.815 ;
        RECT 57.535 121.280 57.785 123.565 ;
        RECT 58.860 123.160 59.190 123.565 ;
        RECT 59.460 123.160 59.790 123.565 ;
        RECT 60.060 123.160 60.390 123.565 ;
        RECT 60.660 123.160 60.990 123.565 ;
        RECT 62.620 123.050 62.850 124.200 ;
        RECT 58.930 122.300 59.390 122.530 ;
        RECT 60.330 122.300 60.790 122.530 ;
        RECT 62.480 122.440 63.080 123.050 ;
        RECT 58.650 121.795 58.880 122.140 ;
        RECT 58.485 121.640 58.880 121.795 ;
        RECT 58.485 121.605 58.865 121.640 ;
        RECT 58.485 121.280 58.675 121.605 ;
        RECT 59.065 121.480 59.255 122.300 ;
        RECT 60.050 121.795 60.280 122.140 ;
        RECT 59.885 121.640 60.280 121.795 ;
        RECT 59.885 121.605 60.265 121.640 ;
        RECT 57.500 120.505 58.675 121.280 ;
        RECT 58.930 121.410 59.390 121.480 ;
        RECT 58.930 121.250 59.415 121.410 ;
        RECT 59.065 121.185 59.415 121.250 ;
        RECT 59.885 121.185 60.075 121.605 ;
        RECT 60.465 121.480 60.655 122.300 ;
        RECT 60.330 121.350 60.790 121.480 ;
        RECT 60.330 121.250 60.810 121.350 ;
        RECT 62.480 121.290 62.675 122.440 ;
        RECT 63.285 122.280 63.475 124.600 ;
        RECT 64.780 124.590 66.115 125.370 ;
        RECT 65.165 124.200 66.115 124.590 ;
        RECT 66.295 125.530 66.610 125.785 ;
        RECT 66.295 124.440 66.485 125.530 ;
        RECT 67.045 125.370 67.235 127.690 ;
        RECT 67.670 127.480 67.900 127.530 ;
        RECT 68.260 127.480 68.490 127.530 ;
        RECT 67.670 127.290 68.490 127.480 ;
        RECT 67.670 125.770 67.900 127.290 ;
        RECT 68.260 125.770 68.490 127.290 ;
        RECT 67.670 125.530 68.490 125.770 ;
        RECT 66.660 124.600 67.620 125.370 ;
        RECT 66.295 124.200 66.610 124.440 ;
        RECT 65.165 122.690 65.355 124.200 ;
        RECT 65.790 122.690 66.020 124.200 ;
        RECT 66.380 123.050 66.610 124.200 ;
        RECT 65.160 122.685 66.100 122.690 ;
        RECT 65.160 122.280 66.105 122.685 ;
        RECT 62.900 122.260 63.860 122.280 ;
        RECT 64.780 122.260 66.105 122.280 ;
        RECT 62.900 122.070 66.105 122.260 ;
        RECT 62.900 122.050 63.860 122.070 ;
        RECT 64.780 122.050 66.105 122.070 ;
        RECT 62.900 121.495 63.860 121.725 ;
        RECT 64.780 121.495 65.740 121.725 ;
        RECT 59.065 120.995 60.075 121.185 ;
        RECT 59.065 120.915 59.415 120.995 ;
        RECT 58.930 120.835 59.415 120.915 ;
        RECT 58.930 120.685 59.390 120.835 ;
        RECT 57.500 120.480 58.860 120.505 ;
        RECT 57.500 120.280 58.880 120.480 ;
        RECT 58.650 119.480 58.880 120.280 ;
        RECT 59.065 119.275 59.255 120.685 ;
        RECT 59.885 120.505 60.075 120.995 ;
        RECT 60.465 121.195 60.810 121.250 ;
        RECT 61.250 121.195 62.250 121.280 ;
        RECT 60.465 121.005 62.250 121.195 ;
        RECT 60.465 120.915 60.810 121.005 ;
        RECT 60.330 120.880 60.810 120.915 ;
        RECT 60.330 120.685 60.790 120.880 ;
        RECT 59.885 120.480 60.265 120.505 ;
        RECT 59.885 120.315 60.280 120.480 ;
        RECT 60.050 119.480 60.280 120.315 ;
        RECT 60.465 119.275 60.655 120.685 ;
        RECT 61.250 120.280 62.250 121.005 ;
        RECT 62.480 120.690 63.080 121.290 ;
        RECT 58.930 119.045 59.390 119.275 ;
        RECT 60.330 119.045 60.790 119.275 ;
        RECT 62.620 117.535 62.850 120.690 ;
        RECT 62.535 117.290 62.850 117.535 ;
        RECT 62.535 116.110 62.725 117.290 ;
        RECT 63.285 117.085 63.475 121.495 ;
        RECT 63.910 121.240 64.140 121.290 ;
        RECT 64.500 121.240 64.730 121.290 ;
        RECT 63.910 121.050 64.730 121.240 ;
        RECT 63.910 117.535 64.140 121.050 ;
        RECT 63.910 117.530 64.255 117.535 ;
        RECT 64.500 117.530 64.730 121.050 ;
        RECT 63.910 117.290 64.730 117.530 ;
        RECT 62.900 116.855 63.860 117.085 ;
        RECT 62.960 116.545 63.800 116.855 ;
        RECT 64.065 116.800 64.605 117.290 ;
        RECT 65.165 117.085 65.355 121.495 ;
        RECT 65.915 121.290 66.105 122.050 ;
        RECT 65.790 121.045 66.105 121.290 ;
        RECT 66.280 122.450 66.890 123.050 ;
        RECT 66.280 122.440 66.610 122.450 ;
        RECT 66.280 121.290 66.470 122.440 ;
        RECT 67.045 122.280 67.235 124.600 ;
        RECT 67.805 124.440 68.365 125.530 ;
        RECT 68.925 125.370 69.115 127.690 ;
        RECT 69.550 125.770 69.780 127.530 ;
        RECT 69.550 125.530 69.865 125.770 ;
        RECT 68.540 124.600 69.500 125.370 ;
        RECT 67.670 124.200 68.490 124.440 ;
        RECT 67.670 122.680 67.900 124.200 ;
        RECT 68.260 122.680 68.490 124.200 ;
        RECT 67.670 122.490 68.490 122.680 ;
        RECT 67.670 122.440 67.900 122.490 ;
        RECT 68.260 122.440 68.490 122.490 ;
        RECT 68.925 122.280 69.115 124.600 ;
        RECT 69.675 124.440 69.865 125.530 ;
        RECT 70.805 125.370 70.995 127.690 ;
        RECT 71.430 125.775 71.660 127.530 ;
        RECT 71.430 125.530 71.745 125.775 ;
        RECT 70.400 124.600 71.400 125.370 ;
        RECT 69.550 124.195 69.865 124.440 ;
        RECT 69.550 122.685 69.780 124.195 ;
        RECT 69.550 122.440 69.875 122.685 ;
        RECT 66.660 122.050 67.620 122.280 ;
        RECT 68.540 122.050 69.500 122.280 ;
        RECT 69.685 121.730 69.875 122.440 ;
        RECT 70.805 122.280 70.995 124.600 ;
        RECT 71.555 124.440 71.745 125.530 ;
        RECT 72.685 125.370 72.875 127.690 ;
        RECT 73.310 125.785 73.540 127.530 ;
        RECT 74.560 127.290 75.420 127.690 ;
        RECT 85.590 127.650 86.490 127.690 ;
        RECT 87.470 127.650 88.660 127.690 ;
        RECT 73.310 125.530 73.625 125.785 ;
        RECT 72.280 124.600 73.280 125.370 ;
        RECT 71.430 124.195 71.745 124.440 ;
        RECT 71.430 123.050 71.660 124.195 ;
        RECT 71.250 122.450 71.850 123.050 ;
        RECT 71.430 122.440 71.660 122.450 ;
        RECT 72.685 122.280 72.875 124.600 ;
        RECT 73.435 124.440 73.625 125.530 ;
        RECT 74.560 125.760 74.755 127.290 ;
        RECT 75.190 125.770 75.420 127.290 ;
        RECT 75.190 125.760 75.515 125.770 ;
        RECT 74.560 125.370 75.515 125.760 ;
        RECT 74.160 124.600 75.515 125.370 ;
        RECT 76.070 125.035 76.720 125.220 ;
        RECT 77.670 125.035 77.990 125.070 ;
        RECT 76.070 124.845 77.990 125.035 ;
        RECT 76.070 124.670 76.720 124.845 ;
        RECT 77.670 124.810 77.990 124.845 ;
        RECT 73.310 124.200 73.625 124.440 ;
        RECT 73.310 123.050 73.540 124.200 ;
        RECT 74.560 124.195 75.515 124.600 ;
        RECT 78.880 124.590 79.230 126.810 ;
        RECT 85.280 125.765 85.510 127.530 ;
        RECT 85.195 125.530 85.510 125.765 ;
        RECT 85.195 124.440 85.385 125.530 ;
        RECT 85.945 125.370 86.135 127.650 ;
        RECT 87.820 127.530 88.660 127.650 ;
        RECT 87.820 127.300 88.680 127.530 ;
        RECT 87.825 125.770 88.015 127.300 ;
        RECT 88.450 125.775 88.680 127.300 ;
        RECT 89.040 125.785 89.270 127.530 ;
        RECT 88.450 125.770 88.775 125.775 ;
        RECT 87.825 125.370 88.775 125.770 ;
        RECT 85.560 124.600 86.520 125.370 ;
        RECT 74.560 124.190 75.510 124.195 ;
        RECT 73.130 122.450 73.730 123.050 ;
        RECT 74.560 122.670 74.755 124.190 ;
        RECT 75.190 122.670 75.420 124.190 ;
        RECT 81.520 123.815 81.850 124.220 ;
        RECT 82.120 123.815 82.450 124.220 ;
        RECT 82.720 123.815 83.050 124.220 ;
        RECT 83.320 123.815 83.650 124.220 ;
        RECT 85.195 124.200 85.510 124.440 ;
        RECT 73.310 122.440 73.540 122.450 ;
        RECT 74.560 122.280 75.420 122.670 ;
        RECT 80.195 123.565 83.650 123.815 ;
        RECT 70.400 122.050 75.420 122.280 ;
        RECT 66.660 121.500 69.875 121.730 ;
        RECT 66.660 121.495 67.620 121.500 ;
        RECT 68.540 121.495 69.875 121.500 ;
        RECT 70.420 121.495 71.380 121.725 ;
        RECT 72.300 121.690 73.260 121.725 ;
        RECT 72.300 121.495 73.510 121.690 ;
        RECT 66.280 121.280 66.610 121.290 ;
        RECT 65.790 117.525 66.020 121.045 ;
        RECT 66.280 120.680 66.890 121.280 ;
        RECT 66.380 117.525 66.610 120.680 ;
        RECT 65.790 117.290 66.105 117.525 ;
        RECT 64.780 116.855 65.740 117.085 ;
        RECT 64.055 116.610 64.605 116.800 ;
        RECT 62.900 116.315 63.860 116.545 ;
        RECT 62.535 115.870 62.850 116.110 ;
        RECT 62.620 112.110 62.850 115.870 ;
        RECT 63.285 111.905 63.475 116.315 ;
        RECT 64.065 116.110 64.605 116.610 ;
        RECT 64.790 116.545 65.730 116.855 ;
        RECT 64.780 116.315 65.740 116.545 ;
        RECT 63.910 115.875 64.730 116.110 ;
        RECT 63.910 115.870 64.255 115.875 ;
        RECT 63.910 112.350 64.140 115.870 ;
        RECT 64.500 112.350 64.730 115.875 ;
        RECT 63.910 112.160 64.730 112.350 ;
        RECT 63.910 112.110 64.140 112.160 ;
        RECT 64.500 112.110 64.730 112.160 ;
        RECT 65.165 111.905 65.355 116.315 ;
        RECT 65.915 116.110 66.105 117.290 ;
        RECT 65.790 115.865 66.105 116.110 ;
        RECT 66.275 117.290 66.610 117.525 ;
        RECT 66.275 116.110 66.465 117.290 ;
        RECT 67.045 117.090 67.235 121.495 ;
        RECT 68.920 121.060 69.875 121.495 ;
        RECT 68.925 117.530 69.115 121.060 ;
        RECT 69.550 121.050 69.875 121.060 ;
        RECT 69.550 117.530 69.780 121.050 ;
        RECT 68.925 117.525 69.860 117.530 ;
        RECT 68.925 117.520 69.865 117.525 ;
        RECT 68.920 117.090 69.865 117.520 ;
        RECT 70.805 117.090 70.995 121.495 ;
        RECT 72.680 121.350 73.510 121.495 ;
        RECT 71.240 120.750 71.850 121.350 ;
        RECT 72.680 121.060 73.730 121.350 ;
        RECT 71.430 117.495 71.660 120.750 ;
        RECT 72.685 117.530 72.875 121.060 ;
        RECT 73.120 120.750 73.730 121.060 ;
        RECT 73.310 117.535 73.540 120.750 ;
        RECT 74.100 119.385 74.350 122.050 ;
        RECT 74.870 119.360 76.060 121.520 ;
        RECT 78.880 120.090 79.230 122.310 ;
        RECT 80.195 121.280 80.445 123.565 ;
        RECT 81.520 123.160 81.850 123.565 ;
        RECT 82.120 123.160 82.450 123.565 ;
        RECT 82.720 123.160 83.050 123.565 ;
        RECT 83.320 123.160 83.650 123.565 ;
        RECT 85.280 123.050 85.510 124.200 ;
        RECT 81.590 122.300 82.050 122.530 ;
        RECT 82.990 122.300 83.450 122.530 ;
        RECT 85.140 122.440 85.740 123.050 ;
        RECT 81.310 121.795 81.540 122.140 ;
        RECT 81.145 121.640 81.540 121.795 ;
        RECT 81.145 121.605 81.525 121.640 ;
        RECT 81.145 121.280 81.335 121.605 ;
        RECT 81.725 121.480 81.915 122.300 ;
        RECT 82.710 121.795 82.940 122.140 ;
        RECT 82.545 121.640 82.940 121.795 ;
        RECT 82.545 121.605 82.925 121.640 ;
        RECT 80.160 120.505 81.335 121.280 ;
        RECT 81.590 121.410 82.050 121.480 ;
        RECT 81.590 121.250 82.075 121.410 ;
        RECT 81.725 121.185 82.075 121.250 ;
        RECT 82.545 121.185 82.735 121.605 ;
        RECT 83.125 121.480 83.315 122.300 ;
        RECT 82.990 121.350 83.450 121.480 ;
        RECT 82.990 121.250 83.470 121.350 ;
        RECT 85.140 121.290 85.335 122.440 ;
        RECT 85.945 122.280 86.135 124.600 ;
        RECT 87.440 124.590 88.775 125.370 ;
        RECT 87.825 124.200 88.775 124.590 ;
        RECT 88.955 125.530 89.270 125.785 ;
        RECT 88.955 124.440 89.145 125.530 ;
        RECT 89.705 125.370 89.895 127.690 ;
        RECT 90.330 127.480 90.560 127.530 ;
        RECT 90.920 127.480 91.150 127.530 ;
        RECT 90.330 127.290 91.150 127.480 ;
        RECT 90.330 125.770 90.560 127.290 ;
        RECT 90.920 125.770 91.150 127.290 ;
        RECT 90.330 125.530 91.150 125.770 ;
        RECT 89.320 124.600 90.280 125.370 ;
        RECT 88.955 124.200 89.270 124.440 ;
        RECT 87.825 122.690 88.015 124.200 ;
        RECT 88.450 122.690 88.680 124.200 ;
        RECT 89.040 123.050 89.270 124.200 ;
        RECT 87.820 122.685 88.760 122.690 ;
        RECT 87.820 122.280 88.765 122.685 ;
        RECT 85.560 122.260 86.520 122.280 ;
        RECT 87.440 122.260 88.765 122.280 ;
        RECT 85.560 122.070 88.765 122.260 ;
        RECT 85.560 122.050 86.520 122.070 ;
        RECT 87.440 122.050 88.765 122.070 ;
        RECT 85.560 121.495 86.520 121.725 ;
        RECT 87.440 121.495 88.400 121.725 ;
        RECT 81.725 120.995 82.735 121.185 ;
        RECT 81.725 120.915 82.075 120.995 ;
        RECT 81.590 120.835 82.075 120.915 ;
        RECT 81.590 120.685 82.050 120.835 ;
        RECT 80.160 120.480 81.520 120.505 ;
        RECT 80.160 120.280 81.540 120.480 ;
        RECT 81.310 119.480 81.540 120.280 ;
        RECT 81.725 119.275 81.915 120.685 ;
        RECT 82.545 120.505 82.735 120.995 ;
        RECT 83.125 121.195 83.470 121.250 ;
        RECT 83.910 121.195 84.910 121.280 ;
        RECT 83.125 121.005 84.910 121.195 ;
        RECT 83.125 120.915 83.470 121.005 ;
        RECT 82.990 120.880 83.470 120.915 ;
        RECT 82.990 120.685 83.450 120.880 ;
        RECT 82.545 120.480 82.925 120.505 ;
        RECT 82.545 120.315 82.940 120.480 ;
        RECT 82.710 119.480 82.940 120.315 ;
        RECT 83.125 119.275 83.315 120.685 ;
        RECT 83.910 120.280 84.910 121.005 ;
        RECT 85.140 120.690 85.740 121.290 ;
        RECT 81.590 119.045 82.050 119.275 ;
        RECT 82.990 119.045 83.450 119.275 ;
        RECT 73.310 117.530 73.625 117.535 ;
        RECT 71.430 117.290 71.745 117.495 ;
        RECT 66.660 116.310 67.620 117.090 ;
        RECT 68.540 116.310 69.865 117.090 ;
        RECT 70.400 116.310 71.400 117.090 ;
        RECT 66.275 115.870 66.610 116.110 ;
        RECT 65.790 112.110 66.020 115.865 ;
        RECT 66.380 112.110 66.610 115.870 ;
        RECT 67.045 111.910 67.235 116.310 ;
        RECT 68.925 115.865 69.865 116.310 ;
        RECT 68.925 115.860 69.860 115.865 ;
        RECT 68.925 112.340 69.115 115.860 ;
        RECT 69.550 112.340 69.780 115.860 ;
        RECT 68.925 112.110 69.780 112.340 ;
        RECT 68.925 111.910 69.750 112.110 ;
        RECT 62.900 111.675 63.860 111.905 ;
        RECT 64.780 111.675 65.740 111.905 ;
        RECT 66.660 111.580 67.620 111.910 ;
        RECT 68.540 111.890 69.750 111.910 ;
        RECT 70.805 111.905 70.995 116.310 ;
        RECT 71.555 116.110 71.745 117.290 ;
        RECT 72.685 117.090 73.625 117.530 ;
        RECT 72.280 116.310 73.625 117.090 ;
        RECT 78.880 116.800 79.230 119.020 ;
        RECT 85.280 117.535 85.510 120.690 ;
        RECT 85.195 117.290 85.510 117.535 ;
        RECT 71.430 115.870 71.745 116.110 ;
        RECT 72.685 115.870 73.625 116.310 ;
        RECT 85.195 116.110 85.385 117.290 ;
        RECT 85.945 117.085 86.135 121.495 ;
        RECT 86.570 121.240 86.800 121.290 ;
        RECT 87.160 121.240 87.390 121.290 ;
        RECT 86.570 121.050 87.390 121.240 ;
        RECT 86.570 117.535 86.800 121.050 ;
        RECT 86.570 117.530 86.915 117.535 ;
        RECT 87.160 117.530 87.390 121.050 ;
        RECT 86.570 117.290 87.390 117.530 ;
        RECT 85.560 116.855 86.520 117.085 ;
        RECT 85.620 116.545 86.460 116.855 ;
        RECT 86.725 116.800 87.265 117.290 ;
        RECT 87.825 117.085 88.015 121.495 ;
        RECT 88.575 121.290 88.765 122.050 ;
        RECT 88.450 121.045 88.765 121.290 ;
        RECT 88.940 122.450 89.550 123.050 ;
        RECT 88.940 122.440 89.270 122.450 ;
        RECT 88.940 121.290 89.130 122.440 ;
        RECT 89.705 122.280 89.895 124.600 ;
        RECT 90.465 124.440 91.025 125.530 ;
        RECT 91.585 125.370 91.775 127.690 ;
        RECT 92.210 125.770 92.440 127.530 ;
        RECT 92.210 125.530 92.525 125.770 ;
        RECT 91.200 124.600 92.160 125.370 ;
        RECT 90.330 124.200 91.150 124.440 ;
        RECT 90.330 122.680 90.560 124.200 ;
        RECT 90.920 122.680 91.150 124.200 ;
        RECT 90.330 122.490 91.150 122.680 ;
        RECT 90.330 122.440 90.560 122.490 ;
        RECT 90.920 122.440 91.150 122.490 ;
        RECT 91.585 122.280 91.775 124.600 ;
        RECT 92.335 124.440 92.525 125.530 ;
        RECT 93.465 125.370 93.655 127.690 ;
        RECT 94.090 125.775 94.320 127.530 ;
        RECT 94.090 125.530 94.405 125.775 ;
        RECT 93.060 124.600 94.060 125.370 ;
        RECT 92.210 124.195 92.525 124.440 ;
        RECT 92.210 122.685 92.440 124.195 ;
        RECT 92.210 122.440 92.535 122.685 ;
        RECT 89.320 122.050 90.280 122.280 ;
        RECT 91.200 122.050 92.160 122.280 ;
        RECT 92.345 121.730 92.535 122.440 ;
        RECT 93.465 122.280 93.655 124.600 ;
        RECT 94.215 124.440 94.405 125.530 ;
        RECT 95.345 125.370 95.535 127.690 ;
        RECT 95.970 125.785 96.200 127.530 ;
        RECT 97.220 127.290 98.080 127.690 ;
        RECT 108.250 127.650 109.150 127.690 ;
        RECT 110.130 127.650 111.320 127.690 ;
        RECT 95.970 125.530 96.285 125.785 ;
        RECT 94.940 124.600 95.940 125.370 ;
        RECT 94.090 124.195 94.405 124.440 ;
        RECT 94.090 123.050 94.320 124.195 ;
        RECT 93.910 122.450 94.510 123.050 ;
        RECT 94.090 122.440 94.320 122.450 ;
        RECT 95.345 122.280 95.535 124.600 ;
        RECT 96.095 124.440 96.285 125.530 ;
        RECT 97.220 125.760 97.415 127.290 ;
        RECT 97.850 125.770 98.080 127.290 ;
        RECT 97.850 125.760 98.175 125.770 ;
        RECT 97.220 125.370 98.175 125.760 ;
        RECT 96.820 124.600 98.175 125.370 ;
        RECT 98.730 125.035 99.380 125.220 ;
        RECT 100.330 125.035 100.650 125.070 ;
        RECT 98.730 124.845 100.650 125.035 ;
        RECT 98.730 124.670 99.380 124.845 ;
        RECT 100.330 124.810 100.650 124.845 ;
        RECT 95.970 124.200 96.285 124.440 ;
        RECT 95.970 123.050 96.200 124.200 ;
        RECT 97.220 124.195 98.175 124.600 ;
        RECT 101.540 124.590 101.890 126.810 ;
        RECT 107.940 125.765 108.170 127.530 ;
        RECT 107.855 125.530 108.170 125.765 ;
        RECT 107.855 124.440 108.045 125.530 ;
        RECT 108.605 125.370 108.795 127.650 ;
        RECT 110.480 127.530 111.320 127.650 ;
        RECT 110.480 127.300 111.340 127.530 ;
        RECT 110.485 125.770 110.675 127.300 ;
        RECT 111.110 125.775 111.340 127.300 ;
        RECT 111.700 125.785 111.930 127.530 ;
        RECT 111.110 125.770 111.435 125.775 ;
        RECT 110.485 125.370 111.435 125.770 ;
        RECT 108.220 124.600 109.180 125.370 ;
        RECT 97.220 124.190 98.170 124.195 ;
        RECT 95.790 122.450 96.390 123.050 ;
        RECT 97.220 122.670 97.415 124.190 ;
        RECT 97.850 122.670 98.080 124.190 ;
        RECT 104.180 123.815 104.510 124.220 ;
        RECT 104.780 123.815 105.110 124.220 ;
        RECT 105.380 123.815 105.710 124.220 ;
        RECT 105.980 123.815 106.310 124.220 ;
        RECT 107.855 124.200 108.170 124.440 ;
        RECT 95.970 122.440 96.200 122.450 ;
        RECT 97.220 122.280 98.080 122.670 ;
        RECT 102.855 123.565 106.310 123.815 ;
        RECT 93.060 122.050 98.080 122.280 ;
        RECT 89.320 121.500 92.535 121.730 ;
        RECT 89.320 121.495 90.280 121.500 ;
        RECT 91.200 121.495 92.535 121.500 ;
        RECT 93.080 121.495 94.040 121.725 ;
        RECT 94.960 121.690 95.920 121.725 ;
        RECT 94.960 121.495 96.170 121.690 ;
        RECT 88.940 121.280 89.270 121.290 ;
        RECT 88.450 117.525 88.680 121.045 ;
        RECT 88.940 120.680 89.550 121.280 ;
        RECT 89.040 117.525 89.270 120.680 ;
        RECT 88.450 117.290 88.765 117.525 ;
        RECT 87.440 116.855 88.400 117.085 ;
        RECT 86.715 116.610 87.265 116.800 ;
        RECT 85.560 116.315 86.520 116.545 ;
        RECT 85.195 115.870 85.510 116.110 ;
        RECT 71.430 112.110 71.660 115.870 ;
        RECT 72.685 112.340 72.875 115.870 ;
        RECT 73.310 115.865 73.625 115.870 ;
        RECT 73.310 112.340 73.540 115.865 ;
        RECT 72.680 111.905 73.540 112.340 ;
        RECT 68.540 111.680 69.630 111.890 ;
        RECT 68.540 111.580 69.500 111.680 ;
        RECT 70.420 111.675 71.380 111.905 ;
        RECT 72.300 111.680 73.540 111.905 ;
        RECT 72.300 111.675 73.260 111.680 ;
        RECT 74.040 111.110 75.230 113.270 ;
        RECT 75.700 111.110 76.890 113.270 ;
        RECT 78.880 112.300 79.230 114.520 ;
        RECT 85.280 112.110 85.510 115.870 ;
        RECT 85.945 111.905 86.135 116.315 ;
        RECT 86.725 116.110 87.265 116.610 ;
        RECT 87.450 116.545 88.390 116.855 ;
        RECT 87.440 116.315 88.400 116.545 ;
        RECT 86.570 115.875 87.390 116.110 ;
        RECT 86.570 115.870 86.915 115.875 ;
        RECT 86.570 112.350 86.800 115.870 ;
        RECT 87.160 112.350 87.390 115.875 ;
        RECT 86.570 112.160 87.390 112.350 ;
        RECT 86.570 112.110 86.800 112.160 ;
        RECT 87.160 112.110 87.390 112.160 ;
        RECT 87.825 111.905 88.015 116.315 ;
        RECT 88.575 116.110 88.765 117.290 ;
        RECT 88.450 115.865 88.765 116.110 ;
        RECT 88.935 117.290 89.270 117.525 ;
        RECT 88.935 116.110 89.125 117.290 ;
        RECT 89.705 117.090 89.895 121.495 ;
        RECT 91.580 121.060 92.535 121.495 ;
        RECT 91.585 117.530 91.775 121.060 ;
        RECT 92.210 121.050 92.535 121.060 ;
        RECT 92.210 117.530 92.440 121.050 ;
        RECT 91.585 117.525 92.520 117.530 ;
        RECT 91.585 117.520 92.525 117.525 ;
        RECT 91.580 117.090 92.525 117.520 ;
        RECT 93.465 117.090 93.655 121.495 ;
        RECT 95.340 121.350 96.170 121.495 ;
        RECT 93.900 120.750 94.510 121.350 ;
        RECT 95.340 121.060 96.390 121.350 ;
        RECT 94.090 117.495 94.320 120.750 ;
        RECT 95.345 117.530 95.535 121.060 ;
        RECT 95.780 120.750 96.390 121.060 ;
        RECT 95.970 117.535 96.200 120.750 ;
        RECT 96.760 119.385 97.010 122.050 ;
        RECT 97.530 119.360 98.720 121.520 ;
        RECT 101.540 120.090 101.890 122.310 ;
        RECT 102.855 121.280 103.105 123.565 ;
        RECT 104.180 123.160 104.510 123.565 ;
        RECT 104.780 123.160 105.110 123.565 ;
        RECT 105.380 123.160 105.710 123.565 ;
        RECT 105.980 123.160 106.310 123.565 ;
        RECT 107.940 123.050 108.170 124.200 ;
        RECT 104.250 122.300 104.710 122.530 ;
        RECT 105.650 122.300 106.110 122.530 ;
        RECT 107.800 122.440 108.400 123.050 ;
        RECT 103.970 121.795 104.200 122.140 ;
        RECT 103.805 121.640 104.200 121.795 ;
        RECT 103.805 121.605 104.185 121.640 ;
        RECT 103.805 121.280 103.995 121.605 ;
        RECT 104.385 121.480 104.575 122.300 ;
        RECT 105.370 121.795 105.600 122.140 ;
        RECT 105.205 121.640 105.600 121.795 ;
        RECT 105.205 121.605 105.585 121.640 ;
        RECT 102.820 120.505 103.995 121.280 ;
        RECT 104.250 121.410 104.710 121.480 ;
        RECT 104.250 121.250 104.735 121.410 ;
        RECT 104.385 121.185 104.735 121.250 ;
        RECT 105.205 121.185 105.395 121.605 ;
        RECT 105.785 121.480 105.975 122.300 ;
        RECT 105.650 121.350 106.110 121.480 ;
        RECT 105.650 121.250 106.130 121.350 ;
        RECT 107.800 121.290 107.995 122.440 ;
        RECT 108.605 122.280 108.795 124.600 ;
        RECT 110.100 124.590 111.435 125.370 ;
        RECT 110.485 124.200 111.435 124.590 ;
        RECT 111.615 125.530 111.930 125.785 ;
        RECT 111.615 124.440 111.805 125.530 ;
        RECT 112.365 125.370 112.555 127.690 ;
        RECT 112.990 127.480 113.220 127.530 ;
        RECT 113.580 127.480 113.810 127.530 ;
        RECT 112.990 127.290 113.810 127.480 ;
        RECT 112.990 125.770 113.220 127.290 ;
        RECT 113.580 125.770 113.810 127.290 ;
        RECT 112.990 125.530 113.810 125.770 ;
        RECT 111.980 124.600 112.940 125.370 ;
        RECT 111.615 124.200 111.930 124.440 ;
        RECT 110.485 122.690 110.675 124.200 ;
        RECT 111.110 122.690 111.340 124.200 ;
        RECT 111.700 123.050 111.930 124.200 ;
        RECT 110.480 122.685 111.420 122.690 ;
        RECT 110.480 122.280 111.425 122.685 ;
        RECT 108.220 122.260 109.180 122.280 ;
        RECT 110.100 122.260 111.425 122.280 ;
        RECT 108.220 122.070 111.425 122.260 ;
        RECT 108.220 122.050 109.180 122.070 ;
        RECT 110.100 122.050 111.425 122.070 ;
        RECT 108.220 121.495 109.180 121.725 ;
        RECT 110.100 121.495 111.060 121.725 ;
        RECT 104.385 120.995 105.395 121.185 ;
        RECT 104.385 120.915 104.735 120.995 ;
        RECT 104.250 120.835 104.735 120.915 ;
        RECT 104.250 120.685 104.710 120.835 ;
        RECT 102.820 120.480 104.180 120.505 ;
        RECT 102.820 120.280 104.200 120.480 ;
        RECT 103.970 119.480 104.200 120.280 ;
        RECT 104.385 119.275 104.575 120.685 ;
        RECT 105.205 120.505 105.395 120.995 ;
        RECT 105.785 121.195 106.130 121.250 ;
        RECT 106.570 121.195 107.570 121.280 ;
        RECT 105.785 121.005 107.570 121.195 ;
        RECT 105.785 120.915 106.130 121.005 ;
        RECT 105.650 120.880 106.130 120.915 ;
        RECT 105.650 120.685 106.110 120.880 ;
        RECT 105.205 120.480 105.585 120.505 ;
        RECT 105.205 120.315 105.600 120.480 ;
        RECT 105.370 119.480 105.600 120.315 ;
        RECT 105.785 119.275 105.975 120.685 ;
        RECT 106.570 120.280 107.570 121.005 ;
        RECT 107.800 120.690 108.400 121.290 ;
        RECT 104.250 119.045 104.710 119.275 ;
        RECT 105.650 119.045 106.110 119.275 ;
        RECT 95.970 117.530 96.285 117.535 ;
        RECT 94.090 117.290 94.405 117.495 ;
        RECT 89.320 116.310 90.280 117.090 ;
        RECT 91.200 116.310 92.525 117.090 ;
        RECT 93.060 116.310 94.060 117.090 ;
        RECT 88.935 115.870 89.270 116.110 ;
        RECT 88.450 112.110 88.680 115.865 ;
        RECT 89.040 112.110 89.270 115.870 ;
        RECT 89.705 111.910 89.895 116.310 ;
        RECT 91.585 115.865 92.525 116.310 ;
        RECT 91.585 115.860 92.520 115.865 ;
        RECT 91.585 112.340 91.775 115.860 ;
        RECT 92.210 112.340 92.440 115.860 ;
        RECT 91.585 112.110 92.440 112.340 ;
        RECT 91.585 111.910 92.410 112.110 ;
        RECT 85.560 111.675 86.520 111.905 ;
        RECT 87.440 111.675 88.400 111.905 ;
        RECT 89.320 111.580 90.280 111.910 ;
        RECT 91.200 111.890 92.410 111.910 ;
        RECT 93.465 111.905 93.655 116.310 ;
        RECT 94.215 116.110 94.405 117.290 ;
        RECT 95.345 117.090 96.285 117.530 ;
        RECT 94.940 116.310 96.285 117.090 ;
        RECT 101.540 116.800 101.890 119.020 ;
        RECT 107.940 117.535 108.170 120.690 ;
        RECT 107.855 117.290 108.170 117.535 ;
        RECT 94.090 115.870 94.405 116.110 ;
        RECT 95.345 115.870 96.285 116.310 ;
        RECT 107.855 116.110 108.045 117.290 ;
        RECT 108.605 117.085 108.795 121.495 ;
        RECT 109.230 121.240 109.460 121.290 ;
        RECT 109.820 121.240 110.050 121.290 ;
        RECT 109.230 121.050 110.050 121.240 ;
        RECT 109.230 117.535 109.460 121.050 ;
        RECT 109.230 117.530 109.575 117.535 ;
        RECT 109.820 117.530 110.050 121.050 ;
        RECT 109.230 117.290 110.050 117.530 ;
        RECT 108.220 116.855 109.180 117.085 ;
        RECT 108.280 116.545 109.120 116.855 ;
        RECT 109.385 116.800 109.925 117.290 ;
        RECT 110.485 117.085 110.675 121.495 ;
        RECT 111.235 121.290 111.425 122.050 ;
        RECT 111.110 121.045 111.425 121.290 ;
        RECT 111.600 122.450 112.210 123.050 ;
        RECT 111.600 122.440 111.930 122.450 ;
        RECT 111.600 121.290 111.790 122.440 ;
        RECT 112.365 122.280 112.555 124.600 ;
        RECT 113.125 124.440 113.685 125.530 ;
        RECT 114.245 125.370 114.435 127.690 ;
        RECT 114.870 125.770 115.100 127.530 ;
        RECT 114.870 125.530 115.185 125.770 ;
        RECT 113.860 124.600 114.820 125.370 ;
        RECT 112.990 124.200 113.810 124.440 ;
        RECT 112.990 122.680 113.220 124.200 ;
        RECT 113.580 122.680 113.810 124.200 ;
        RECT 112.990 122.490 113.810 122.680 ;
        RECT 112.990 122.440 113.220 122.490 ;
        RECT 113.580 122.440 113.810 122.490 ;
        RECT 114.245 122.280 114.435 124.600 ;
        RECT 114.995 124.440 115.185 125.530 ;
        RECT 116.125 125.370 116.315 127.690 ;
        RECT 116.750 125.775 116.980 127.530 ;
        RECT 116.750 125.530 117.065 125.775 ;
        RECT 115.720 124.600 116.720 125.370 ;
        RECT 114.870 124.195 115.185 124.440 ;
        RECT 114.870 122.685 115.100 124.195 ;
        RECT 114.870 122.440 115.195 122.685 ;
        RECT 111.980 122.050 112.940 122.280 ;
        RECT 113.860 122.050 114.820 122.280 ;
        RECT 115.005 121.730 115.195 122.440 ;
        RECT 116.125 122.280 116.315 124.600 ;
        RECT 116.875 124.440 117.065 125.530 ;
        RECT 118.005 125.370 118.195 127.690 ;
        RECT 118.630 125.785 118.860 127.530 ;
        RECT 119.880 127.290 120.740 127.690 ;
        RECT 118.630 125.530 118.945 125.785 ;
        RECT 117.600 124.600 118.600 125.370 ;
        RECT 116.750 124.195 117.065 124.440 ;
        RECT 116.750 123.050 116.980 124.195 ;
        RECT 116.570 122.450 117.170 123.050 ;
        RECT 116.750 122.440 116.980 122.450 ;
        RECT 118.005 122.280 118.195 124.600 ;
        RECT 118.755 124.440 118.945 125.530 ;
        RECT 119.880 125.760 120.075 127.290 ;
        RECT 120.510 125.770 120.740 127.290 ;
        RECT 120.510 125.760 120.835 125.770 ;
        RECT 119.880 125.370 120.835 125.760 ;
        RECT 119.480 124.600 120.835 125.370 ;
        RECT 121.390 125.035 122.040 125.220 ;
        RECT 122.990 125.035 123.310 125.070 ;
        RECT 121.390 124.845 123.310 125.035 ;
        RECT 121.390 124.670 122.040 124.845 ;
        RECT 122.990 124.810 123.310 124.845 ;
        RECT 118.630 124.200 118.945 124.440 ;
        RECT 118.630 123.050 118.860 124.200 ;
        RECT 119.880 124.195 120.835 124.600 ;
        RECT 119.880 124.190 120.830 124.195 ;
        RECT 118.450 122.450 119.050 123.050 ;
        RECT 119.880 122.670 120.075 124.190 ;
        RECT 120.510 122.670 120.740 124.190 ;
        RECT 118.630 122.440 118.860 122.450 ;
        RECT 119.880 122.280 120.740 122.670 ;
        RECT 115.720 122.050 120.740 122.280 ;
        RECT 111.980 121.500 115.195 121.730 ;
        RECT 111.980 121.495 112.940 121.500 ;
        RECT 113.860 121.495 115.195 121.500 ;
        RECT 115.740 121.495 116.700 121.725 ;
        RECT 117.620 121.690 118.580 121.725 ;
        RECT 117.620 121.495 118.830 121.690 ;
        RECT 111.600 121.280 111.930 121.290 ;
        RECT 111.110 117.525 111.340 121.045 ;
        RECT 111.600 120.680 112.210 121.280 ;
        RECT 111.700 117.525 111.930 120.680 ;
        RECT 111.110 117.290 111.425 117.525 ;
        RECT 110.100 116.855 111.060 117.085 ;
        RECT 109.375 116.610 109.925 116.800 ;
        RECT 108.220 116.315 109.180 116.545 ;
        RECT 107.855 115.870 108.170 116.110 ;
        RECT 94.090 112.110 94.320 115.870 ;
        RECT 95.345 112.340 95.535 115.870 ;
        RECT 95.970 115.865 96.285 115.870 ;
        RECT 95.970 112.340 96.200 115.865 ;
        RECT 95.340 111.905 96.200 112.340 ;
        RECT 91.200 111.680 92.290 111.890 ;
        RECT 91.200 111.580 92.160 111.680 ;
        RECT 93.080 111.675 94.040 111.905 ;
        RECT 94.960 111.680 96.200 111.905 ;
        RECT 94.960 111.675 95.920 111.680 ;
        RECT 96.700 111.110 97.890 113.270 ;
        RECT 98.360 111.110 99.550 113.270 ;
        RECT 101.540 112.300 101.890 114.520 ;
        RECT 107.940 112.110 108.170 115.870 ;
        RECT 108.605 111.905 108.795 116.315 ;
        RECT 109.385 116.110 109.925 116.610 ;
        RECT 110.110 116.545 111.050 116.855 ;
        RECT 110.100 116.315 111.060 116.545 ;
        RECT 109.230 115.875 110.050 116.110 ;
        RECT 109.230 115.870 109.575 115.875 ;
        RECT 109.230 112.350 109.460 115.870 ;
        RECT 109.820 112.350 110.050 115.875 ;
        RECT 109.230 112.160 110.050 112.350 ;
        RECT 109.230 112.110 109.460 112.160 ;
        RECT 109.820 112.110 110.050 112.160 ;
        RECT 110.485 111.905 110.675 116.315 ;
        RECT 111.235 116.110 111.425 117.290 ;
        RECT 111.110 115.865 111.425 116.110 ;
        RECT 111.595 117.290 111.930 117.525 ;
        RECT 111.595 116.110 111.785 117.290 ;
        RECT 112.365 117.090 112.555 121.495 ;
        RECT 114.240 121.060 115.195 121.495 ;
        RECT 114.245 117.530 114.435 121.060 ;
        RECT 114.870 121.050 115.195 121.060 ;
        RECT 114.870 117.530 115.100 121.050 ;
        RECT 114.245 117.525 115.180 117.530 ;
        RECT 114.245 117.520 115.185 117.525 ;
        RECT 114.240 117.090 115.185 117.520 ;
        RECT 116.125 117.090 116.315 121.495 ;
        RECT 118.000 121.350 118.830 121.495 ;
        RECT 116.560 120.750 117.170 121.350 ;
        RECT 118.000 121.060 119.050 121.350 ;
        RECT 116.750 117.495 116.980 120.750 ;
        RECT 118.005 117.530 118.195 121.060 ;
        RECT 118.440 120.750 119.050 121.060 ;
        RECT 118.630 117.535 118.860 120.750 ;
        RECT 119.420 119.385 119.670 122.050 ;
        RECT 120.190 119.360 121.380 121.520 ;
        RECT 124.200 120.090 124.550 122.310 ;
        RECT 118.630 117.530 118.945 117.535 ;
        RECT 116.750 117.290 117.065 117.495 ;
        RECT 111.980 116.310 112.940 117.090 ;
        RECT 113.860 116.310 115.185 117.090 ;
        RECT 115.720 116.310 116.720 117.090 ;
        RECT 111.595 115.870 111.930 116.110 ;
        RECT 111.110 112.110 111.340 115.865 ;
        RECT 111.700 112.110 111.930 115.870 ;
        RECT 112.365 111.910 112.555 116.310 ;
        RECT 114.245 115.865 115.185 116.310 ;
        RECT 114.245 115.860 115.180 115.865 ;
        RECT 114.245 112.340 114.435 115.860 ;
        RECT 114.870 112.340 115.100 115.860 ;
        RECT 114.245 112.110 115.100 112.340 ;
        RECT 114.245 111.910 115.070 112.110 ;
        RECT 108.220 111.675 109.180 111.905 ;
        RECT 110.100 111.675 111.060 111.905 ;
        RECT 111.980 111.580 112.940 111.910 ;
        RECT 113.860 111.890 115.070 111.910 ;
        RECT 116.125 111.905 116.315 116.310 ;
        RECT 116.875 116.110 117.065 117.290 ;
        RECT 118.005 117.090 118.945 117.530 ;
        RECT 117.600 116.310 118.945 117.090 ;
        RECT 124.200 116.800 124.550 119.020 ;
        RECT 116.750 115.870 117.065 116.110 ;
        RECT 118.005 115.870 118.945 116.310 ;
        RECT 116.750 112.110 116.980 115.870 ;
        RECT 118.005 112.340 118.195 115.870 ;
        RECT 118.630 115.865 118.945 115.870 ;
        RECT 118.630 112.340 118.860 115.865 ;
        RECT 118.000 111.905 118.860 112.340 ;
        RECT 113.860 111.680 114.950 111.890 ;
        RECT 113.860 111.580 114.820 111.680 ;
        RECT 115.740 111.675 116.700 111.905 ;
        RECT 117.620 111.680 118.860 111.905 ;
        RECT 117.620 111.675 118.580 111.680 ;
        RECT 119.360 111.110 120.550 113.270 ;
        RECT 121.020 111.110 122.210 113.270 ;
        RECT 124.200 112.300 124.550 114.520 ;
        RECT 40.270 110.580 41.170 110.630 ;
        RECT 42.150 110.580 43.050 110.630 ;
        RECT 40.240 110.350 41.200 110.580 ;
        RECT 42.120 110.555 43.080 110.580 ;
        RECT 42.120 110.350 43.340 110.555 ;
        RECT 44.000 110.350 44.960 110.580 ;
        RECT 45.880 110.350 46.840 110.580 ;
        RECT 47.740 110.350 48.740 110.670 ;
        RECT 49.620 110.350 50.620 110.670 ;
        RECT 51.500 110.580 52.500 110.670 ;
        RECT 62.930 110.580 63.830 110.630 ;
        RECT 64.810 110.580 65.710 110.630 ;
        RECT 51.500 110.350 52.760 110.580 ;
        RECT 62.900 110.350 63.860 110.580 ;
        RECT 64.780 110.555 65.740 110.580 ;
        RECT 64.780 110.350 66.000 110.555 ;
        RECT 66.660 110.350 67.620 110.580 ;
        RECT 68.540 110.350 69.500 110.580 ;
        RECT 70.400 110.350 71.400 110.670 ;
        RECT 72.280 110.350 73.280 110.670 ;
        RECT 74.160 110.580 75.160 110.670 ;
        RECT 85.590 110.580 86.490 110.630 ;
        RECT 87.470 110.580 88.370 110.630 ;
        RECT 74.160 110.350 75.420 110.580 ;
        RECT 85.560 110.350 86.520 110.580 ;
        RECT 87.440 110.555 88.400 110.580 ;
        RECT 87.440 110.350 88.660 110.555 ;
        RECT 89.320 110.350 90.280 110.580 ;
        RECT 91.200 110.350 92.160 110.580 ;
        RECT 93.060 110.350 94.060 110.670 ;
        RECT 94.940 110.350 95.940 110.670 ;
        RECT 96.820 110.580 97.820 110.670 ;
        RECT 108.250 110.580 109.150 110.630 ;
        RECT 110.130 110.580 111.030 110.630 ;
        RECT 96.820 110.350 98.080 110.580 ;
        RECT 108.220 110.350 109.180 110.580 ;
        RECT 110.100 110.555 111.060 110.580 ;
        RECT 110.100 110.350 111.320 110.555 ;
        RECT 111.980 110.350 112.940 110.580 ;
        RECT 113.860 110.350 114.820 110.580 ;
        RECT 115.720 110.350 116.720 110.670 ;
        RECT 117.600 110.350 118.600 110.670 ;
        RECT 119.480 110.580 120.480 110.670 ;
        RECT 119.480 110.350 120.740 110.580 ;
        RECT 40.270 110.310 41.170 110.350 ;
        RECT 42.150 110.310 43.340 110.350 ;
        RECT 39.960 108.425 40.190 110.190 ;
        RECT 39.875 108.190 40.190 108.425 ;
        RECT 39.875 107.100 40.065 108.190 ;
        RECT 40.625 108.030 40.815 110.310 ;
        RECT 42.500 110.190 43.340 110.310 ;
        RECT 42.500 109.960 43.360 110.190 ;
        RECT 42.505 108.430 42.695 109.960 ;
        RECT 43.130 108.435 43.360 109.960 ;
        RECT 43.720 108.445 43.950 110.190 ;
        RECT 43.130 108.430 43.455 108.435 ;
        RECT 42.505 108.030 43.455 108.430 ;
        RECT 40.240 107.260 41.200 108.030 ;
        RECT 36.200 106.475 36.530 106.880 ;
        RECT 36.800 106.475 37.130 106.880 ;
        RECT 37.400 106.475 37.730 106.880 ;
        RECT 38.000 106.475 38.330 106.880 ;
        RECT 39.875 106.860 40.190 107.100 ;
        RECT 34.875 106.225 38.330 106.475 ;
        RECT 34.875 103.940 35.125 106.225 ;
        RECT 36.200 105.820 36.530 106.225 ;
        RECT 36.800 105.820 37.130 106.225 ;
        RECT 37.400 105.820 37.730 106.225 ;
        RECT 38.000 105.820 38.330 106.225 ;
        RECT 39.960 105.710 40.190 106.860 ;
        RECT 36.270 104.960 36.730 105.190 ;
        RECT 37.670 104.960 38.130 105.190 ;
        RECT 39.820 105.100 40.420 105.710 ;
        RECT 35.990 104.455 36.220 104.800 ;
        RECT 35.825 104.300 36.220 104.455 ;
        RECT 35.825 104.265 36.205 104.300 ;
        RECT 35.825 103.940 36.015 104.265 ;
        RECT 36.405 104.140 36.595 104.960 ;
        RECT 37.390 104.455 37.620 104.800 ;
        RECT 37.225 104.300 37.620 104.455 ;
        RECT 37.225 104.265 37.605 104.300 ;
        RECT 34.840 103.165 36.015 103.940 ;
        RECT 36.270 104.070 36.730 104.140 ;
        RECT 36.270 103.910 36.755 104.070 ;
        RECT 36.405 103.845 36.755 103.910 ;
        RECT 37.225 103.845 37.415 104.265 ;
        RECT 37.805 104.140 37.995 104.960 ;
        RECT 37.670 104.010 38.130 104.140 ;
        RECT 37.670 103.910 38.150 104.010 ;
        RECT 39.820 103.950 40.015 105.100 ;
        RECT 40.625 104.940 40.815 107.260 ;
        RECT 42.120 107.250 43.455 108.030 ;
        RECT 42.505 106.860 43.455 107.250 ;
        RECT 43.635 108.190 43.950 108.445 ;
        RECT 43.635 107.100 43.825 108.190 ;
        RECT 44.385 108.030 44.575 110.350 ;
        RECT 45.010 110.140 45.240 110.190 ;
        RECT 45.600 110.140 45.830 110.190 ;
        RECT 45.010 109.950 45.830 110.140 ;
        RECT 45.010 108.430 45.240 109.950 ;
        RECT 45.600 108.430 45.830 109.950 ;
        RECT 45.010 108.190 45.830 108.430 ;
        RECT 44.000 107.260 44.960 108.030 ;
        RECT 43.635 106.860 43.950 107.100 ;
        RECT 42.505 105.350 42.695 106.860 ;
        RECT 43.130 105.350 43.360 106.860 ;
        RECT 43.720 105.710 43.950 106.860 ;
        RECT 42.500 105.345 43.440 105.350 ;
        RECT 42.500 104.940 43.445 105.345 ;
        RECT 40.240 104.920 41.200 104.940 ;
        RECT 42.120 104.920 43.445 104.940 ;
        RECT 40.240 104.730 43.445 104.920 ;
        RECT 40.240 104.710 41.200 104.730 ;
        RECT 42.120 104.710 43.445 104.730 ;
        RECT 40.240 104.155 41.200 104.385 ;
        RECT 42.120 104.155 43.080 104.385 ;
        RECT 36.405 103.655 37.415 103.845 ;
        RECT 36.405 103.575 36.755 103.655 ;
        RECT 36.270 103.495 36.755 103.575 ;
        RECT 36.270 103.345 36.730 103.495 ;
        RECT 34.840 103.140 36.200 103.165 ;
        RECT 34.840 102.940 36.220 103.140 ;
        RECT 35.990 102.140 36.220 102.940 ;
        RECT 36.405 101.935 36.595 103.345 ;
        RECT 37.225 103.165 37.415 103.655 ;
        RECT 37.805 103.855 38.150 103.910 ;
        RECT 38.590 103.855 39.590 103.940 ;
        RECT 37.805 103.665 39.590 103.855 ;
        RECT 37.805 103.575 38.150 103.665 ;
        RECT 37.670 103.540 38.150 103.575 ;
        RECT 37.670 103.345 38.130 103.540 ;
        RECT 37.225 103.140 37.605 103.165 ;
        RECT 37.225 102.975 37.620 103.140 ;
        RECT 37.390 102.140 37.620 102.975 ;
        RECT 37.805 101.935 37.995 103.345 ;
        RECT 38.590 102.940 39.590 103.665 ;
        RECT 39.820 103.350 40.420 103.950 ;
        RECT 36.270 101.705 36.730 101.935 ;
        RECT 37.670 101.705 38.130 101.935 ;
        RECT 39.960 100.195 40.190 103.350 ;
        RECT 39.875 99.950 40.190 100.195 ;
        RECT 39.875 98.770 40.065 99.950 ;
        RECT 40.625 99.745 40.815 104.155 ;
        RECT 41.250 103.900 41.480 103.950 ;
        RECT 41.840 103.900 42.070 103.950 ;
        RECT 41.250 103.710 42.070 103.900 ;
        RECT 41.250 100.195 41.480 103.710 ;
        RECT 41.250 100.190 41.595 100.195 ;
        RECT 41.840 100.190 42.070 103.710 ;
        RECT 41.250 99.950 42.070 100.190 ;
        RECT 40.240 99.515 41.200 99.745 ;
        RECT 40.300 99.205 41.140 99.515 ;
        RECT 41.405 99.460 41.945 99.950 ;
        RECT 42.505 99.745 42.695 104.155 ;
        RECT 43.255 103.950 43.445 104.710 ;
        RECT 43.130 103.705 43.445 103.950 ;
        RECT 43.620 105.110 44.230 105.710 ;
        RECT 43.620 105.100 43.950 105.110 ;
        RECT 43.620 103.950 43.810 105.100 ;
        RECT 44.385 104.940 44.575 107.260 ;
        RECT 45.145 107.100 45.705 108.190 ;
        RECT 46.265 108.030 46.455 110.350 ;
        RECT 46.890 108.430 47.120 110.190 ;
        RECT 46.890 108.190 47.205 108.430 ;
        RECT 45.880 107.260 46.840 108.030 ;
        RECT 45.010 106.860 45.830 107.100 ;
        RECT 45.010 105.340 45.240 106.860 ;
        RECT 45.600 105.340 45.830 106.860 ;
        RECT 45.010 105.150 45.830 105.340 ;
        RECT 45.010 105.100 45.240 105.150 ;
        RECT 45.600 105.100 45.830 105.150 ;
        RECT 46.265 104.940 46.455 107.260 ;
        RECT 47.015 107.100 47.205 108.190 ;
        RECT 48.145 108.030 48.335 110.350 ;
        RECT 48.770 108.435 49.000 110.190 ;
        RECT 48.770 108.190 49.085 108.435 ;
        RECT 47.740 107.260 48.740 108.030 ;
        RECT 46.890 106.855 47.205 107.100 ;
        RECT 46.890 105.345 47.120 106.855 ;
        RECT 46.890 105.100 47.215 105.345 ;
        RECT 44.000 104.710 44.960 104.940 ;
        RECT 45.880 104.710 46.840 104.940 ;
        RECT 47.025 104.390 47.215 105.100 ;
        RECT 48.145 104.940 48.335 107.260 ;
        RECT 48.895 107.100 49.085 108.190 ;
        RECT 50.025 108.030 50.215 110.350 ;
        RECT 50.650 108.445 50.880 110.190 ;
        RECT 51.900 109.950 52.760 110.350 ;
        RECT 62.930 110.310 63.830 110.350 ;
        RECT 64.810 110.310 66.000 110.350 ;
        RECT 50.650 108.190 50.965 108.445 ;
        RECT 49.620 107.260 50.620 108.030 ;
        RECT 48.770 106.855 49.085 107.100 ;
        RECT 48.770 105.710 49.000 106.855 ;
        RECT 48.590 105.110 49.190 105.710 ;
        RECT 48.770 105.100 49.000 105.110 ;
        RECT 50.025 104.940 50.215 107.260 ;
        RECT 50.775 107.100 50.965 108.190 ;
        RECT 51.900 108.420 52.095 109.950 ;
        RECT 52.530 108.430 52.760 109.950 ;
        RECT 52.530 108.420 52.855 108.430 ;
        RECT 62.620 108.425 62.850 110.190 ;
        RECT 51.900 108.030 52.855 108.420 ;
        RECT 51.500 107.260 52.855 108.030 ;
        RECT 62.535 108.190 62.850 108.425 ;
        RECT 53.410 107.695 54.060 107.880 ;
        RECT 55.010 107.695 55.330 107.730 ;
        RECT 53.410 107.505 55.330 107.695 ;
        RECT 53.410 107.330 54.060 107.505 ;
        RECT 55.010 107.470 55.330 107.505 ;
        RECT 50.650 106.860 50.965 107.100 ;
        RECT 50.650 105.710 50.880 106.860 ;
        RECT 51.900 106.855 52.855 107.260 ;
        RECT 62.535 107.100 62.725 108.190 ;
        RECT 63.285 108.030 63.475 110.310 ;
        RECT 65.160 110.190 66.000 110.310 ;
        RECT 65.160 109.960 66.020 110.190 ;
        RECT 65.165 108.430 65.355 109.960 ;
        RECT 65.790 108.435 66.020 109.960 ;
        RECT 66.380 108.445 66.610 110.190 ;
        RECT 65.790 108.430 66.115 108.435 ;
        RECT 65.165 108.030 66.115 108.430 ;
        RECT 62.900 107.260 63.860 108.030 ;
        RECT 51.900 106.850 52.850 106.855 ;
        RECT 50.470 105.110 51.070 105.710 ;
        RECT 51.900 105.330 52.095 106.850 ;
        RECT 52.530 105.330 52.760 106.850 ;
        RECT 58.860 106.475 59.190 106.880 ;
        RECT 59.460 106.475 59.790 106.880 ;
        RECT 60.060 106.475 60.390 106.880 ;
        RECT 60.660 106.475 60.990 106.880 ;
        RECT 62.535 106.860 62.850 107.100 ;
        RECT 50.650 105.100 50.880 105.110 ;
        RECT 51.900 104.940 52.760 105.330 ;
        RECT 57.535 106.225 60.990 106.475 ;
        RECT 47.740 104.710 52.760 104.940 ;
        RECT 44.000 104.160 47.215 104.390 ;
        RECT 44.000 104.155 44.960 104.160 ;
        RECT 45.880 104.155 47.215 104.160 ;
        RECT 47.760 104.155 48.720 104.385 ;
        RECT 49.640 104.350 50.600 104.385 ;
        RECT 49.640 104.155 50.850 104.350 ;
        RECT 43.620 103.940 43.950 103.950 ;
        RECT 43.130 100.185 43.360 103.705 ;
        RECT 43.620 103.340 44.230 103.940 ;
        RECT 43.720 100.185 43.950 103.340 ;
        RECT 43.130 99.950 43.445 100.185 ;
        RECT 42.120 99.515 43.080 99.745 ;
        RECT 41.395 99.270 41.945 99.460 ;
        RECT 40.240 98.975 41.200 99.205 ;
        RECT 39.875 98.530 40.190 98.770 ;
        RECT 39.960 94.770 40.190 98.530 ;
        RECT 40.625 94.565 40.815 98.975 ;
        RECT 41.405 98.770 41.945 99.270 ;
        RECT 42.130 99.205 43.070 99.515 ;
        RECT 42.120 98.975 43.080 99.205 ;
        RECT 41.250 98.535 42.070 98.770 ;
        RECT 41.250 98.530 41.595 98.535 ;
        RECT 41.250 95.010 41.480 98.530 ;
        RECT 41.840 95.010 42.070 98.535 ;
        RECT 41.250 94.820 42.070 95.010 ;
        RECT 41.250 94.770 41.480 94.820 ;
        RECT 41.840 94.770 42.070 94.820 ;
        RECT 42.505 94.565 42.695 98.975 ;
        RECT 43.255 98.770 43.445 99.950 ;
        RECT 43.130 98.525 43.445 98.770 ;
        RECT 43.615 99.950 43.950 100.185 ;
        RECT 43.615 98.770 43.805 99.950 ;
        RECT 44.385 99.750 44.575 104.155 ;
        RECT 46.260 103.720 47.215 104.155 ;
        RECT 46.265 100.190 46.455 103.720 ;
        RECT 46.890 103.710 47.215 103.720 ;
        RECT 46.890 100.190 47.120 103.710 ;
        RECT 46.265 100.185 47.200 100.190 ;
        RECT 46.265 100.180 47.205 100.185 ;
        RECT 46.260 99.750 47.205 100.180 ;
        RECT 48.145 99.750 48.335 104.155 ;
        RECT 50.020 104.010 50.850 104.155 ;
        RECT 48.580 103.410 49.190 104.010 ;
        RECT 50.020 103.720 51.070 104.010 ;
        RECT 48.770 100.155 49.000 103.410 ;
        RECT 50.025 100.190 50.215 103.720 ;
        RECT 50.460 103.410 51.070 103.720 ;
        RECT 50.650 100.195 50.880 103.410 ;
        RECT 51.440 102.045 51.690 104.710 ;
        RECT 52.210 102.020 53.400 104.180 ;
        RECT 56.220 102.750 56.570 104.970 ;
        RECT 57.535 103.940 57.785 106.225 ;
        RECT 58.860 105.820 59.190 106.225 ;
        RECT 59.460 105.820 59.790 106.225 ;
        RECT 60.060 105.820 60.390 106.225 ;
        RECT 60.660 105.820 60.990 106.225 ;
        RECT 62.620 105.710 62.850 106.860 ;
        RECT 58.930 104.960 59.390 105.190 ;
        RECT 60.330 104.960 60.790 105.190 ;
        RECT 62.480 105.100 63.080 105.710 ;
        RECT 58.650 104.455 58.880 104.800 ;
        RECT 58.485 104.300 58.880 104.455 ;
        RECT 58.485 104.265 58.865 104.300 ;
        RECT 58.485 103.940 58.675 104.265 ;
        RECT 59.065 104.140 59.255 104.960 ;
        RECT 60.050 104.455 60.280 104.800 ;
        RECT 59.885 104.300 60.280 104.455 ;
        RECT 59.885 104.265 60.265 104.300 ;
        RECT 57.500 103.165 58.675 103.940 ;
        RECT 58.930 104.070 59.390 104.140 ;
        RECT 58.930 103.910 59.415 104.070 ;
        RECT 59.065 103.845 59.415 103.910 ;
        RECT 59.885 103.845 60.075 104.265 ;
        RECT 60.465 104.140 60.655 104.960 ;
        RECT 60.330 104.010 60.790 104.140 ;
        RECT 60.330 103.910 60.810 104.010 ;
        RECT 62.480 103.950 62.675 105.100 ;
        RECT 63.285 104.940 63.475 107.260 ;
        RECT 64.780 107.250 66.115 108.030 ;
        RECT 65.165 106.860 66.115 107.250 ;
        RECT 66.295 108.190 66.610 108.445 ;
        RECT 66.295 107.100 66.485 108.190 ;
        RECT 67.045 108.030 67.235 110.350 ;
        RECT 67.670 110.140 67.900 110.190 ;
        RECT 68.260 110.140 68.490 110.190 ;
        RECT 67.670 109.950 68.490 110.140 ;
        RECT 67.670 108.430 67.900 109.950 ;
        RECT 68.260 108.430 68.490 109.950 ;
        RECT 67.670 108.190 68.490 108.430 ;
        RECT 66.660 107.260 67.620 108.030 ;
        RECT 66.295 106.860 66.610 107.100 ;
        RECT 65.165 105.350 65.355 106.860 ;
        RECT 65.790 105.350 66.020 106.860 ;
        RECT 66.380 105.710 66.610 106.860 ;
        RECT 65.160 105.345 66.100 105.350 ;
        RECT 65.160 104.940 66.105 105.345 ;
        RECT 62.900 104.920 63.860 104.940 ;
        RECT 64.780 104.920 66.105 104.940 ;
        RECT 62.900 104.730 66.105 104.920 ;
        RECT 62.900 104.710 63.860 104.730 ;
        RECT 64.780 104.710 66.105 104.730 ;
        RECT 62.900 104.155 63.860 104.385 ;
        RECT 64.780 104.155 65.740 104.385 ;
        RECT 59.065 103.655 60.075 103.845 ;
        RECT 59.065 103.575 59.415 103.655 ;
        RECT 58.930 103.495 59.415 103.575 ;
        RECT 58.930 103.345 59.390 103.495 ;
        RECT 57.500 103.140 58.860 103.165 ;
        RECT 57.500 102.940 58.880 103.140 ;
        RECT 58.650 102.140 58.880 102.940 ;
        RECT 59.065 101.935 59.255 103.345 ;
        RECT 59.885 103.165 60.075 103.655 ;
        RECT 60.465 103.855 60.810 103.910 ;
        RECT 61.250 103.855 62.250 103.940 ;
        RECT 60.465 103.665 62.250 103.855 ;
        RECT 60.465 103.575 60.810 103.665 ;
        RECT 60.330 103.540 60.810 103.575 ;
        RECT 60.330 103.345 60.790 103.540 ;
        RECT 59.885 103.140 60.265 103.165 ;
        RECT 59.885 102.975 60.280 103.140 ;
        RECT 60.050 102.140 60.280 102.975 ;
        RECT 60.465 101.935 60.655 103.345 ;
        RECT 61.250 102.940 62.250 103.665 ;
        RECT 62.480 103.350 63.080 103.950 ;
        RECT 58.930 101.705 59.390 101.935 ;
        RECT 60.330 101.705 60.790 101.935 ;
        RECT 50.650 100.190 50.965 100.195 ;
        RECT 48.770 99.950 49.085 100.155 ;
        RECT 44.000 98.970 44.960 99.750 ;
        RECT 45.880 98.970 47.205 99.750 ;
        RECT 47.740 98.970 48.740 99.750 ;
        RECT 43.615 98.530 43.950 98.770 ;
        RECT 43.130 94.770 43.360 98.525 ;
        RECT 43.720 94.770 43.950 98.530 ;
        RECT 44.385 94.570 44.575 98.970 ;
        RECT 46.265 98.525 47.205 98.970 ;
        RECT 46.265 98.520 47.200 98.525 ;
        RECT 46.265 95.000 46.455 98.520 ;
        RECT 46.890 95.000 47.120 98.520 ;
        RECT 46.265 94.770 47.120 95.000 ;
        RECT 46.265 94.570 47.090 94.770 ;
        RECT 40.240 94.335 41.200 94.565 ;
        RECT 42.120 94.335 43.080 94.565 ;
        RECT 44.000 94.240 44.960 94.570 ;
        RECT 45.880 94.550 47.090 94.570 ;
        RECT 48.145 94.565 48.335 98.970 ;
        RECT 48.895 98.770 49.085 99.950 ;
        RECT 50.025 99.750 50.965 100.190 ;
        RECT 49.620 98.970 50.965 99.750 ;
        RECT 56.220 99.460 56.570 101.680 ;
        RECT 62.620 100.195 62.850 103.350 ;
        RECT 62.535 99.950 62.850 100.195 ;
        RECT 48.770 98.530 49.085 98.770 ;
        RECT 50.025 98.530 50.965 98.970 ;
        RECT 62.535 98.770 62.725 99.950 ;
        RECT 63.285 99.745 63.475 104.155 ;
        RECT 63.910 103.900 64.140 103.950 ;
        RECT 64.500 103.900 64.730 103.950 ;
        RECT 63.910 103.710 64.730 103.900 ;
        RECT 63.910 100.195 64.140 103.710 ;
        RECT 63.910 100.190 64.255 100.195 ;
        RECT 64.500 100.190 64.730 103.710 ;
        RECT 63.910 99.950 64.730 100.190 ;
        RECT 62.900 99.515 63.860 99.745 ;
        RECT 62.960 99.205 63.800 99.515 ;
        RECT 64.065 99.460 64.605 99.950 ;
        RECT 65.165 99.745 65.355 104.155 ;
        RECT 65.915 103.950 66.105 104.710 ;
        RECT 65.790 103.705 66.105 103.950 ;
        RECT 66.280 105.110 66.890 105.710 ;
        RECT 66.280 105.100 66.610 105.110 ;
        RECT 66.280 103.950 66.470 105.100 ;
        RECT 67.045 104.940 67.235 107.260 ;
        RECT 67.805 107.100 68.365 108.190 ;
        RECT 68.925 108.030 69.115 110.350 ;
        RECT 69.550 108.430 69.780 110.190 ;
        RECT 69.550 108.190 69.865 108.430 ;
        RECT 68.540 107.260 69.500 108.030 ;
        RECT 67.670 106.860 68.490 107.100 ;
        RECT 67.670 105.340 67.900 106.860 ;
        RECT 68.260 105.340 68.490 106.860 ;
        RECT 67.670 105.150 68.490 105.340 ;
        RECT 67.670 105.100 67.900 105.150 ;
        RECT 68.260 105.100 68.490 105.150 ;
        RECT 68.925 104.940 69.115 107.260 ;
        RECT 69.675 107.100 69.865 108.190 ;
        RECT 70.805 108.030 70.995 110.350 ;
        RECT 71.430 108.435 71.660 110.190 ;
        RECT 71.430 108.190 71.745 108.435 ;
        RECT 70.400 107.260 71.400 108.030 ;
        RECT 69.550 106.855 69.865 107.100 ;
        RECT 69.550 105.345 69.780 106.855 ;
        RECT 69.550 105.100 69.875 105.345 ;
        RECT 66.660 104.710 67.620 104.940 ;
        RECT 68.540 104.710 69.500 104.940 ;
        RECT 69.685 104.390 69.875 105.100 ;
        RECT 70.805 104.940 70.995 107.260 ;
        RECT 71.555 107.100 71.745 108.190 ;
        RECT 72.685 108.030 72.875 110.350 ;
        RECT 73.310 108.445 73.540 110.190 ;
        RECT 74.560 109.950 75.420 110.350 ;
        RECT 85.590 110.310 86.490 110.350 ;
        RECT 87.470 110.310 88.660 110.350 ;
        RECT 73.310 108.190 73.625 108.445 ;
        RECT 72.280 107.260 73.280 108.030 ;
        RECT 71.430 106.855 71.745 107.100 ;
        RECT 71.430 105.710 71.660 106.855 ;
        RECT 71.250 105.110 71.850 105.710 ;
        RECT 71.430 105.100 71.660 105.110 ;
        RECT 72.685 104.940 72.875 107.260 ;
        RECT 73.435 107.100 73.625 108.190 ;
        RECT 74.560 108.420 74.755 109.950 ;
        RECT 75.190 108.430 75.420 109.950 ;
        RECT 75.190 108.420 75.515 108.430 ;
        RECT 74.560 108.030 75.515 108.420 ;
        RECT 74.160 107.260 75.515 108.030 ;
        RECT 76.070 107.695 76.720 107.880 ;
        RECT 77.670 107.695 77.990 107.730 ;
        RECT 76.070 107.505 77.990 107.695 ;
        RECT 76.070 107.330 76.720 107.505 ;
        RECT 77.670 107.470 77.990 107.505 ;
        RECT 73.310 106.860 73.625 107.100 ;
        RECT 73.310 105.710 73.540 106.860 ;
        RECT 74.560 106.855 75.515 107.260 ;
        RECT 78.880 107.250 79.230 109.470 ;
        RECT 85.280 108.425 85.510 110.190 ;
        RECT 85.195 108.190 85.510 108.425 ;
        RECT 85.195 107.100 85.385 108.190 ;
        RECT 85.945 108.030 86.135 110.310 ;
        RECT 87.820 110.190 88.660 110.310 ;
        RECT 87.820 109.960 88.680 110.190 ;
        RECT 87.825 108.430 88.015 109.960 ;
        RECT 88.450 108.435 88.680 109.960 ;
        RECT 89.040 108.445 89.270 110.190 ;
        RECT 88.450 108.430 88.775 108.435 ;
        RECT 87.825 108.030 88.775 108.430 ;
        RECT 85.560 107.260 86.520 108.030 ;
        RECT 74.560 106.850 75.510 106.855 ;
        RECT 73.130 105.110 73.730 105.710 ;
        RECT 74.560 105.330 74.755 106.850 ;
        RECT 75.190 105.330 75.420 106.850 ;
        RECT 81.520 106.475 81.850 106.880 ;
        RECT 82.120 106.475 82.450 106.880 ;
        RECT 82.720 106.475 83.050 106.880 ;
        RECT 83.320 106.475 83.650 106.880 ;
        RECT 85.195 106.860 85.510 107.100 ;
        RECT 73.310 105.100 73.540 105.110 ;
        RECT 74.560 104.940 75.420 105.330 ;
        RECT 80.195 106.225 83.650 106.475 ;
        RECT 70.400 104.710 75.420 104.940 ;
        RECT 66.660 104.160 69.875 104.390 ;
        RECT 66.660 104.155 67.620 104.160 ;
        RECT 68.540 104.155 69.875 104.160 ;
        RECT 70.420 104.155 71.380 104.385 ;
        RECT 72.300 104.350 73.260 104.385 ;
        RECT 72.300 104.155 73.510 104.350 ;
        RECT 66.280 103.940 66.610 103.950 ;
        RECT 65.790 100.185 66.020 103.705 ;
        RECT 66.280 103.340 66.890 103.940 ;
        RECT 66.380 100.185 66.610 103.340 ;
        RECT 65.790 99.950 66.105 100.185 ;
        RECT 64.780 99.515 65.740 99.745 ;
        RECT 64.055 99.270 64.605 99.460 ;
        RECT 62.900 98.975 63.860 99.205 ;
        RECT 62.535 98.530 62.850 98.770 ;
        RECT 48.770 94.770 49.000 98.530 ;
        RECT 50.025 95.000 50.215 98.530 ;
        RECT 50.650 98.525 50.965 98.530 ;
        RECT 50.650 95.000 50.880 98.525 ;
        RECT 50.020 94.565 50.880 95.000 ;
        RECT 45.880 94.340 46.970 94.550 ;
        RECT 45.880 94.240 46.840 94.340 ;
        RECT 47.760 94.335 48.720 94.565 ;
        RECT 49.640 94.340 50.880 94.565 ;
        RECT 49.640 94.335 50.600 94.340 ;
        RECT 51.380 93.770 52.570 95.930 ;
        RECT 53.040 93.770 54.230 95.930 ;
        RECT 56.220 94.960 56.570 97.180 ;
        RECT 62.620 94.770 62.850 98.530 ;
        RECT 63.285 94.565 63.475 98.975 ;
        RECT 64.065 98.770 64.605 99.270 ;
        RECT 64.790 99.205 65.730 99.515 ;
        RECT 64.780 98.975 65.740 99.205 ;
        RECT 63.910 98.535 64.730 98.770 ;
        RECT 63.910 98.530 64.255 98.535 ;
        RECT 63.910 95.010 64.140 98.530 ;
        RECT 64.500 95.010 64.730 98.535 ;
        RECT 63.910 94.820 64.730 95.010 ;
        RECT 63.910 94.770 64.140 94.820 ;
        RECT 64.500 94.770 64.730 94.820 ;
        RECT 65.165 94.565 65.355 98.975 ;
        RECT 65.915 98.770 66.105 99.950 ;
        RECT 65.790 98.525 66.105 98.770 ;
        RECT 66.275 99.950 66.610 100.185 ;
        RECT 66.275 98.770 66.465 99.950 ;
        RECT 67.045 99.750 67.235 104.155 ;
        RECT 68.920 103.720 69.875 104.155 ;
        RECT 68.925 100.190 69.115 103.720 ;
        RECT 69.550 103.710 69.875 103.720 ;
        RECT 69.550 100.190 69.780 103.710 ;
        RECT 68.925 100.185 69.860 100.190 ;
        RECT 68.925 100.180 69.865 100.185 ;
        RECT 68.920 99.750 69.865 100.180 ;
        RECT 70.805 99.750 70.995 104.155 ;
        RECT 72.680 104.010 73.510 104.155 ;
        RECT 71.240 103.410 71.850 104.010 ;
        RECT 72.680 103.720 73.730 104.010 ;
        RECT 71.430 100.155 71.660 103.410 ;
        RECT 72.685 100.190 72.875 103.720 ;
        RECT 73.120 103.410 73.730 103.720 ;
        RECT 73.310 100.195 73.540 103.410 ;
        RECT 74.100 102.045 74.350 104.710 ;
        RECT 74.870 102.020 76.060 104.180 ;
        RECT 78.880 102.750 79.230 104.970 ;
        RECT 80.195 103.940 80.445 106.225 ;
        RECT 81.520 105.820 81.850 106.225 ;
        RECT 82.120 105.820 82.450 106.225 ;
        RECT 82.720 105.820 83.050 106.225 ;
        RECT 83.320 105.820 83.650 106.225 ;
        RECT 85.280 105.710 85.510 106.860 ;
        RECT 81.590 104.960 82.050 105.190 ;
        RECT 82.990 104.960 83.450 105.190 ;
        RECT 85.140 105.100 85.740 105.710 ;
        RECT 81.310 104.455 81.540 104.800 ;
        RECT 81.145 104.300 81.540 104.455 ;
        RECT 81.145 104.265 81.525 104.300 ;
        RECT 81.145 103.940 81.335 104.265 ;
        RECT 81.725 104.140 81.915 104.960 ;
        RECT 82.710 104.455 82.940 104.800 ;
        RECT 82.545 104.300 82.940 104.455 ;
        RECT 82.545 104.265 82.925 104.300 ;
        RECT 80.160 103.165 81.335 103.940 ;
        RECT 81.590 104.070 82.050 104.140 ;
        RECT 81.590 103.910 82.075 104.070 ;
        RECT 81.725 103.845 82.075 103.910 ;
        RECT 82.545 103.845 82.735 104.265 ;
        RECT 83.125 104.140 83.315 104.960 ;
        RECT 82.990 104.010 83.450 104.140 ;
        RECT 82.990 103.910 83.470 104.010 ;
        RECT 85.140 103.950 85.335 105.100 ;
        RECT 85.945 104.940 86.135 107.260 ;
        RECT 87.440 107.250 88.775 108.030 ;
        RECT 87.825 106.860 88.775 107.250 ;
        RECT 88.955 108.190 89.270 108.445 ;
        RECT 88.955 107.100 89.145 108.190 ;
        RECT 89.705 108.030 89.895 110.350 ;
        RECT 90.330 110.140 90.560 110.190 ;
        RECT 90.920 110.140 91.150 110.190 ;
        RECT 90.330 109.950 91.150 110.140 ;
        RECT 90.330 108.430 90.560 109.950 ;
        RECT 90.920 108.430 91.150 109.950 ;
        RECT 90.330 108.190 91.150 108.430 ;
        RECT 89.320 107.260 90.280 108.030 ;
        RECT 88.955 106.860 89.270 107.100 ;
        RECT 87.825 105.350 88.015 106.860 ;
        RECT 88.450 105.350 88.680 106.860 ;
        RECT 89.040 105.710 89.270 106.860 ;
        RECT 87.820 105.345 88.760 105.350 ;
        RECT 87.820 104.940 88.765 105.345 ;
        RECT 85.560 104.920 86.520 104.940 ;
        RECT 87.440 104.920 88.765 104.940 ;
        RECT 85.560 104.730 88.765 104.920 ;
        RECT 85.560 104.710 86.520 104.730 ;
        RECT 87.440 104.710 88.765 104.730 ;
        RECT 85.560 104.155 86.520 104.385 ;
        RECT 87.440 104.155 88.400 104.385 ;
        RECT 81.725 103.655 82.735 103.845 ;
        RECT 81.725 103.575 82.075 103.655 ;
        RECT 81.590 103.495 82.075 103.575 ;
        RECT 81.590 103.345 82.050 103.495 ;
        RECT 80.160 103.140 81.520 103.165 ;
        RECT 80.160 102.940 81.540 103.140 ;
        RECT 81.310 102.140 81.540 102.940 ;
        RECT 81.725 101.935 81.915 103.345 ;
        RECT 82.545 103.165 82.735 103.655 ;
        RECT 83.125 103.855 83.470 103.910 ;
        RECT 83.910 103.855 84.910 103.940 ;
        RECT 83.125 103.665 84.910 103.855 ;
        RECT 83.125 103.575 83.470 103.665 ;
        RECT 82.990 103.540 83.470 103.575 ;
        RECT 82.990 103.345 83.450 103.540 ;
        RECT 82.545 103.140 82.925 103.165 ;
        RECT 82.545 102.975 82.940 103.140 ;
        RECT 82.710 102.140 82.940 102.975 ;
        RECT 83.125 101.935 83.315 103.345 ;
        RECT 83.910 102.940 84.910 103.665 ;
        RECT 85.140 103.350 85.740 103.950 ;
        RECT 81.590 101.705 82.050 101.935 ;
        RECT 82.990 101.705 83.450 101.935 ;
        RECT 73.310 100.190 73.625 100.195 ;
        RECT 71.430 99.950 71.745 100.155 ;
        RECT 66.660 98.970 67.620 99.750 ;
        RECT 68.540 98.970 69.865 99.750 ;
        RECT 70.400 98.970 71.400 99.750 ;
        RECT 66.275 98.530 66.610 98.770 ;
        RECT 65.790 94.770 66.020 98.525 ;
        RECT 66.380 94.770 66.610 98.530 ;
        RECT 67.045 94.570 67.235 98.970 ;
        RECT 68.925 98.525 69.865 98.970 ;
        RECT 68.925 98.520 69.860 98.525 ;
        RECT 68.925 95.000 69.115 98.520 ;
        RECT 69.550 95.000 69.780 98.520 ;
        RECT 68.925 94.770 69.780 95.000 ;
        RECT 68.925 94.570 69.750 94.770 ;
        RECT 62.900 94.335 63.860 94.565 ;
        RECT 64.780 94.335 65.740 94.565 ;
        RECT 66.660 94.240 67.620 94.570 ;
        RECT 68.540 94.550 69.750 94.570 ;
        RECT 70.805 94.565 70.995 98.970 ;
        RECT 71.555 98.770 71.745 99.950 ;
        RECT 72.685 99.750 73.625 100.190 ;
        RECT 72.280 98.970 73.625 99.750 ;
        RECT 78.880 99.460 79.230 101.680 ;
        RECT 85.280 100.195 85.510 103.350 ;
        RECT 85.195 99.950 85.510 100.195 ;
        RECT 71.430 98.530 71.745 98.770 ;
        RECT 72.685 98.530 73.625 98.970 ;
        RECT 85.195 98.770 85.385 99.950 ;
        RECT 85.945 99.745 86.135 104.155 ;
        RECT 86.570 103.900 86.800 103.950 ;
        RECT 87.160 103.900 87.390 103.950 ;
        RECT 86.570 103.710 87.390 103.900 ;
        RECT 86.570 100.195 86.800 103.710 ;
        RECT 86.570 100.190 86.915 100.195 ;
        RECT 87.160 100.190 87.390 103.710 ;
        RECT 86.570 99.950 87.390 100.190 ;
        RECT 85.560 99.515 86.520 99.745 ;
        RECT 85.620 99.205 86.460 99.515 ;
        RECT 86.725 99.460 87.265 99.950 ;
        RECT 87.825 99.745 88.015 104.155 ;
        RECT 88.575 103.950 88.765 104.710 ;
        RECT 88.450 103.705 88.765 103.950 ;
        RECT 88.940 105.110 89.550 105.710 ;
        RECT 88.940 105.100 89.270 105.110 ;
        RECT 88.940 103.950 89.130 105.100 ;
        RECT 89.705 104.940 89.895 107.260 ;
        RECT 90.465 107.100 91.025 108.190 ;
        RECT 91.585 108.030 91.775 110.350 ;
        RECT 92.210 108.430 92.440 110.190 ;
        RECT 92.210 108.190 92.525 108.430 ;
        RECT 91.200 107.260 92.160 108.030 ;
        RECT 90.330 106.860 91.150 107.100 ;
        RECT 90.330 105.340 90.560 106.860 ;
        RECT 90.920 105.340 91.150 106.860 ;
        RECT 90.330 105.150 91.150 105.340 ;
        RECT 90.330 105.100 90.560 105.150 ;
        RECT 90.920 105.100 91.150 105.150 ;
        RECT 91.585 104.940 91.775 107.260 ;
        RECT 92.335 107.100 92.525 108.190 ;
        RECT 93.465 108.030 93.655 110.350 ;
        RECT 94.090 108.435 94.320 110.190 ;
        RECT 94.090 108.190 94.405 108.435 ;
        RECT 93.060 107.260 94.060 108.030 ;
        RECT 92.210 106.855 92.525 107.100 ;
        RECT 92.210 105.345 92.440 106.855 ;
        RECT 92.210 105.100 92.535 105.345 ;
        RECT 89.320 104.710 90.280 104.940 ;
        RECT 91.200 104.710 92.160 104.940 ;
        RECT 92.345 104.390 92.535 105.100 ;
        RECT 93.465 104.940 93.655 107.260 ;
        RECT 94.215 107.100 94.405 108.190 ;
        RECT 95.345 108.030 95.535 110.350 ;
        RECT 95.970 108.445 96.200 110.190 ;
        RECT 97.220 109.950 98.080 110.350 ;
        RECT 108.250 110.310 109.150 110.350 ;
        RECT 110.130 110.310 111.320 110.350 ;
        RECT 95.970 108.190 96.285 108.445 ;
        RECT 94.940 107.260 95.940 108.030 ;
        RECT 94.090 106.855 94.405 107.100 ;
        RECT 94.090 105.710 94.320 106.855 ;
        RECT 93.910 105.110 94.510 105.710 ;
        RECT 94.090 105.100 94.320 105.110 ;
        RECT 95.345 104.940 95.535 107.260 ;
        RECT 96.095 107.100 96.285 108.190 ;
        RECT 97.220 108.420 97.415 109.950 ;
        RECT 97.850 108.430 98.080 109.950 ;
        RECT 97.850 108.420 98.175 108.430 ;
        RECT 97.220 108.030 98.175 108.420 ;
        RECT 96.820 107.260 98.175 108.030 ;
        RECT 98.730 107.695 99.380 107.880 ;
        RECT 100.330 107.695 100.650 107.730 ;
        RECT 98.730 107.505 100.650 107.695 ;
        RECT 98.730 107.330 99.380 107.505 ;
        RECT 100.330 107.470 100.650 107.505 ;
        RECT 95.970 106.860 96.285 107.100 ;
        RECT 95.970 105.710 96.200 106.860 ;
        RECT 97.220 106.855 98.175 107.260 ;
        RECT 101.540 107.250 101.890 109.470 ;
        RECT 107.940 108.425 108.170 110.190 ;
        RECT 107.855 108.190 108.170 108.425 ;
        RECT 107.855 107.100 108.045 108.190 ;
        RECT 108.605 108.030 108.795 110.310 ;
        RECT 110.480 110.190 111.320 110.310 ;
        RECT 110.480 109.960 111.340 110.190 ;
        RECT 110.485 108.430 110.675 109.960 ;
        RECT 111.110 108.435 111.340 109.960 ;
        RECT 111.700 108.445 111.930 110.190 ;
        RECT 111.110 108.430 111.435 108.435 ;
        RECT 110.485 108.030 111.435 108.430 ;
        RECT 108.220 107.260 109.180 108.030 ;
        RECT 97.220 106.850 98.170 106.855 ;
        RECT 95.790 105.110 96.390 105.710 ;
        RECT 97.220 105.330 97.415 106.850 ;
        RECT 97.850 105.330 98.080 106.850 ;
        RECT 104.180 106.475 104.510 106.880 ;
        RECT 104.780 106.475 105.110 106.880 ;
        RECT 105.380 106.475 105.710 106.880 ;
        RECT 105.980 106.475 106.310 106.880 ;
        RECT 107.855 106.860 108.170 107.100 ;
        RECT 95.970 105.100 96.200 105.110 ;
        RECT 97.220 104.940 98.080 105.330 ;
        RECT 102.855 106.225 106.310 106.475 ;
        RECT 93.060 104.710 98.080 104.940 ;
        RECT 89.320 104.160 92.535 104.390 ;
        RECT 89.320 104.155 90.280 104.160 ;
        RECT 91.200 104.155 92.535 104.160 ;
        RECT 93.080 104.155 94.040 104.385 ;
        RECT 94.960 104.350 95.920 104.385 ;
        RECT 94.960 104.155 96.170 104.350 ;
        RECT 88.940 103.940 89.270 103.950 ;
        RECT 88.450 100.185 88.680 103.705 ;
        RECT 88.940 103.340 89.550 103.940 ;
        RECT 89.040 100.185 89.270 103.340 ;
        RECT 88.450 99.950 88.765 100.185 ;
        RECT 87.440 99.515 88.400 99.745 ;
        RECT 86.715 99.270 87.265 99.460 ;
        RECT 85.560 98.975 86.520 99.205 ;
        RECT 85.195 98.530 85.510 98.770 ;
        RECT 71.430 94.770 71.660 98.530 ;
        RECT 72.685 95.000 72.875 98.530 ;
        RECT 73.310 98.525 73.625 98.530 ;
        RECT 73.310 95.000 73.540 98.525 ;
        RECT 72.680 94.565 73.540 95.000 ;
        RECT 68.540 94.340 69.630 94.550 ;
        RECT 68.540 94.240 69.500 94.340 ;
        RECT 70.420 94.335 71.380 94.565 ;
        RECT 72.300 94.340 73.540 94.565 ;
        RECT 72.300 94.335 73.260 94.340 ;
        RECT 74.040 93.770 75.230 95.930 ;
        RECT 75.700 93.770 76.890 95.930 ;
        RECT 78.880 94.960 79.230 97.180 ;
        RECT 85.280 94.770 85.510 98.530 ;
        RECT 85.945 94.565 86.135 98.975 ;
        RECT 86.725 98.770 87.265 99.270 ;
        RECT 87.450 99.205 88.390 99.515 ;
        RECT 87.440 98.975 88.400 99.205 ;
        RECT 86.570 98.535 87.390 98.770 ;
        RECT 86.570 98.530 86.915 98.535 ;
        RECT 86.570 95.010 86.800 98.530 ;
        RECT 87.160 95.010 87.390 98.535 ;
        RECT 86.570 94.820 87.390 95.010 ;
        RECT 86.570 94.770 86.800 94.820 ;
        RECT 87.160 94.770 87.390 94.820 ;
        RECT 87.825 94.565 88.015 98.975 ;
        RECT 88.575 98.770 88.765 99.950 ;
        RECT 88.450 98.525 88.765 98.770 ;
        RECT 88.935 99.950 89.270 100.185 ;
        RECT 88.935 98.770 89.125 99.950 ;
        RECT 89.705 99.750 89.895 104.155 ;
        RECT 91.580 103.720 92.535 104.155 ;
        RECT 91.585 100.190 91.775 103.720 ;
        RECT 92.210 103.710 92.535 103.720 ;
        RECT 92.210 100.190 92.440 103.710 ;
        RECT 91.585 100.185 92.520 100.190 ;
        RECT 91.585 100.180 92.525 100.185 ;
        RECT 91.580 99.750 92.525 100.180 ;
        RECT 93.465 99.750 93.655 104.155 ;
        RECT 95.340 104.010 96.170 104.155 ;
        RECT 93.900 103.410 94.510 104.010 ;
        RECT 95.340 103.720 96.390 104.010 ;
        RECT 94.090 100.155 94.320 103.410 ;
        RECT 95.345 100.190 95.535 103.720 ;
        RECT 95.780 103.410 96.390 103.720 ;
        RECT 95.970 100.195 96.200 103.410 ;
        RECT 96.760 102.045 97.010 104.710 ;
        RECT 97.530 102.020 98.720 104.180 ;
        RECT 101.540 102.750 101.890 104.970 ;
        RECT 102.855 103.940 103.105 106.225 ;
        RECT 104.180 105.820 104.510 106.225 ;
        RECT 104.780 105.820 105.110 106.225 ;
        RECT 105.380 105.820 105.710 106.225 ;
        RECT 105.980 105.820 106.310 106.225 ;
        RECT 107.940 105.710 108.170 106.860 ;
        RECT 104.250 104.960 104.710 105.190 ;
        RECT 105.650 104.960 106.110 105.190 ;
        RECT 107.800 105.100 108.400 105.710 ;
        RECT 103.970 104.455 104.200 104.800 ;
        RECT 103.805 104.300 104.200 104.455 ;
        RECT 103.805 104.265 104.185 104.300 ;
        RECT 103.805 103.940 103.995 104.265 ;
        RECT 104.385 104.140 104.575 104.960 ;
        RECT 105.370 104.455 105.600 104.800 ;
        RECT 105.205 104.300 105.600 104.455 ;
        RECT 105.205 104.265 105.585 104.300 ;
        RECT 102.820 103.165 103.995 103.940 ;
        RECT 104.250 104.070 104.710 104.140 ;
        RECT 104.250 103.910 104.735 104.070 ;
        RECT 104.385 103.845 104.735 103.910 ;
        RECT 105.205 103.845 105.395 104.265 ;
        RECT 105.785 104.140 105.975 104.960 ;
        RECT 105.650 104.010 106.110 104.140 ;
        RECT 105.650 103.910 106.130 104.010 ;
        RECT 107.800 103.950 107.995 105.100 ;
        RECT 108.605 104.940 108.795 107.260 ;
        RECT 110.100 107.250 111.435 108.030 ;
        RECT 110.485 106.860 111.435 107.250 ;
        RECT 111.615 108.190 111.930 108.445 ;
        RECT 111.615 107.100 111.805 108.190 ;
        RECT 112.365 108.030 112.555 110.350 ;
        RECT 112.990 110.140 113.220 110.190 ;
        RECT 113.580 110.140 113.810 110.190 ;
        RECT 112.990 109.950 113.810 110.140 ;
        RECT 112.990 108.430 113.220 109.950 ;
        RECT 113.580 108.430 113.810 109.950 ;
        RECT 112.990 108.190 113.810 108.430 ;
        RECT 111.980 107.260 112.940 108.030 ;
        RECT 111.615 106.860 111.930 107.100 ;
        RECT 110.485 105.350 110.675 106.860 ;
        RECT 111.110 105.350 111.340 106.860 ;
        RECT 111.700 105.710 111.930 106.860 ;
        RECT 110.480 105.345 111.420 105.350 ;
        RECT 110.480 104.940 111.425 105.345 ;
        RECT 108.220 104.920 109.180 104.940 ;
        RECT 110.100 104.920 111.425 104.940 ;
        RECT 108.220 104.730 111.425 104.920 ;
        RECT 108.220 104.710 109.180 104.730 ;
        RECT 110.100 104.710 111.425 104.730 ;
        RECT 108.220 104.155 109.180 104.385 ;
        RECT 110.100 104.155 111.060 104.385 ;
        RECT 104.385 103.655 105.395 103.845 ;
        RECT 104.385 103.575 104.735 103.655 ;
        RECT 104.250 103.495 104.735 103.575 ;
        RECT 104.250 103.345 104.710 103.495 ;
        RECT 102.820 103.140 104.180 103.165 ;
        RECT 102.820 102.940 104.200 103.140 ;
        RECT 103.970 102.140 104.200 102.940 ;
        RECT 104.385 101.935 104.575 103.345 ;
        RECT 105.205 103.165 105.395 103.655 ;
        RECT 105.785 103.855 106.130 103.910 ;
        RECT 106.570 103.855 107.570 103.940 ;
        RECT 105.785 103.665 107.570 103.855 ;
        RECT 105.785 103.575 106.130 103.665 ;
        RECT 105.650 103.540 106.130 103.575 ;
        RECT 105.650 103.345 106.110 103.540 ;
        RECT 105.205 103.140 105.585 103.165 ;
        RECT 105.205 102.975 105.600 103.140 ;
        RECT 105.370 102.140 105.600 102.975 ;
        RECT 105.785 101.935 105.975 103.345 ;
        RECT 106.570 102.940 107.570 103.665 ;
        RECT 107.800 103.350 108.400 103.950 ;
        RECT 104.250 101.705 104.710 101.935 ;
        RECT 105.650 101.705 106.110 101.935 ;
        RECT 95.970 100.190 96.285 100.195 ;
        RECT 94.090 99.950 94.405 100.155 ;
        RECT 89.320 98.970 90.280 99.750 ;
        RECT 91.200 98.970 92.525 99.750 ;
        RECT 93.060 98.970 94.060 99.750 ;
        RECT 88.935 98.530 89.270 98.770 ;
        RECT 88.450 94.770 88.680 98.525 ;
        RECT 89.040 94.770 89.270 98.530 ;
        RECT 89.705 94.570 89.895 98.970 ;
        RECT 91.585 98.525 92.525 98.970 ;
        RECT 91.585 98.520 92.520 98.525 ;
        RECT 91.585 95.000 91.775 98.520 ;
        RECT 92.210 95.000 92.440 98.520 ;
        RECT 91.585 94.770 92.440 95.000 ;
        RECT 91.585 94.570 92.410 94.770 ;
        RECT 85.560 94.335 86.520 94.565 ;
        RECT 87.440 94.335 88.400 94.565 ;
        RECT 89.320 94.240 90.280 94.570 ;
        RECT 91.200 94.550 92.410 94.570 ;
        RECT 93.465 94.565 93.655 98.970 ;
        RECT 94.215 98.770 94.405 99.950 ;
        RECT 95.345 99.750 96.285 100.190 ;
        RECT 94.940 98.970 96.285 99.750 ;
        RECT 101.540 99.460 101.890 101.680 ;
        RECT 107.940 100.195 108.170 103.350 ;
        RECT 107.855 99.950 108.170 100.195 ;
        RECT 94.090 98.530 94.405 98.770 ;
        RECT 95.345 98.530 96.285 98.970 ;
        RECT 107.855 98.770 108.045 99.950 ;
        RECT 108.605 99.745 108.795 104.155 ;
        RECT 109.230 103.900 109.460 103.950 ;
        RECT 109.820 103.900 110.050 103.950 ;
        RECT 109.230 103.710 110.050 103.900 ;
        RECT 109.230 100.195 109.460 103.710 ;
        RECT 109.230 100.190 109.575 100.195 ;
        RECT 109.820 100.190 110.050 103.710 ;
        RECT 109.230 99.950 110.050 100.190 ;
        RECT 108.220 99.515 109.180 99.745 ;
        RECT 108.280 99.205 109.120 99.515 ;
        RECT 109.385 99.460 109.925 99.950 ;
        RECT 110.485 99.745 110.675 104.155 ;
        RECT 111.235 103.950 111.425 104.710 ;
        RECT 111.110 103.705 111.425 103.950 ;
        RECT 111.600 105.110 112.210 105.710 ;
        RECT 111.600 105.100 111.930 105.110 ;
        RECT 111.600 103.950 111.790 105.100 ;
        RECT 112.365 104.940 112.555 107.260 ;
        RECT 113.125 107.100 113.685 108.190 ;
        RECT 114.245 108.030 114.435 110.350 ;
        RECT 114.870 108.430 115.100 110.190 ;
        RECT 114.870 108.190 115.185 108.430 ;
        RECT 113.860 107.260 114.820 108.030 ;
        RECT 112.990 106.860 113.810 107.100 ;
        RECT 112.990 105.340 113.220 106.860 ;
        RECT 113.580 105.340 113.810 106.860 ;
        RECT 112.990 105.150 113.810 105.340 ;
        RECT 112.990 105.100 113.220 105.150 ;
        RECT 113.580 105.100 113.810 105.150 ;
        RECT 114.245 104.940 114.435 107.260 ;
        RECT 114.995 107.100 115.185 108.190 ;
        RECT 116.125 108.030 116.315 110.350 ;
        RECT 116.750 108.435 116.980 110.190 ;
        RECT 116.750 108.190 117.065 108.435 ;
        RECT 115.720 107.260 116.720 108.030 ;
        RECT 114.870 106.855 115.185 107.100 ;
        RECT 114.870 105.345 115.100 106.855 ;
        RECT 114.870 105.100 115.195 105.345 ;
        RECT 111.980 104.710 112.940 104.940 ;
        RECT 113.860 104.710 114.820 104.940 ;
        RECT 115.005 104.390 115.195 105.100 ;
        RECT 116.125 104.940 116.315 107.260 ;
        RECT 116.875 107.100 117.065 108.190 ;
        RECT 118.005 108.030 118.195 110.350 ;
        RECT 118.630 108.445 118.860 110.190 ;
        RECT 119.880 109.950 120.740 110.350 ;
        RECT 118.630 108.190 118.945 108.445 ;
        RECT 117.600 107.260 118.600 108.030 ;
        RECT 116.750 106.855 117.065 107.100 ;
        RECT 116.750 105.710 116.980 106.855 ;
        RECT 116.570 105.110 117.170 105.710 ;
        RECT 116.750 105.100 116.980 105.110 ;
        RECT 118.005 104.940 118.195 107.260 ;
        RECT 118.755 107.100 118.945 108.190 ;
        RECT 119.880 108.420 120.075 109.950 ;
        RECT 120.510 108.430 120.740 109.950 ;
        RECT 120.510 108.420 120.835 108.430 ;
        RECT 119.880 108.030 120.835 108.420 ;
        RECT 119.480 107.260 120.835 108.030 ;
        RECT 121.390 107.695 122.040 107.880 ;
        RECT 122.990 107.695 123.310 107.730 ;
        RECT 121.390 107.505 123.310 107.695 ;
        RECT 121.390 107.330 122.040 107.505 ;
        RECT 122.990 107.470 123.310 107.505 ;
        RECT 118.630 106.860 118.945 107.100 ;
        RECT 118.630 105.710 118.860 106.860 ;
        RECT 119.880 106.855 120.835 107.260 ;
        RECT 124.200 107.250 124.550 109.470 ;
        RECT 119.880 106.850 120.830 106.855 ;
        RECT 118.450 105.110 119.050 105.710 ;
        RECT 119.880 105.330 120.075 106.850 ;
        RECT 120.510 105.330 120.740 106.850 ;
        RECT 118.630 105.100 118.860 105.110 ;
        RECT 119.880 104.940 120.740 105.330 ;
        RECT 115.720 104.710 120.740 104.940 ;
        RECT 111.980 104.160 115.195 104.390 ;
        RECT 111.980 104.155 112.940 104.160 ;
        RECT 113.860 104.155 115.195 104.160 ;
        RECT 115.740 104.155 116.700 104.385 ;
        RECT 117.620 104.350 118.580 104.385 ;
        RECT 117.620 104.155 118.830 104.350 ;
        RECT 111.600 103.940 111.930 103.950 ;
        RECT 111.110 100.185 111.340 103.705 ;
        RECT 111.600 103.340 112.210 103.940 ;
        RECT 111.700 100.185 111.930 103.340 ;
        RECT 111.110 99.950 111.425 100.185 ;
        RECT 110.100 99.515 111.060 99.745 ;
        RECT 109.375 99.270 109.925 99.460 ;
        RECT 108.220 98.975 109.180 99.205 ;
        RECT 107.855 98.530 108.170 98.770 ;
        RECT 94.090 94.770 94.320 98.530 ;
        RECT 95.345 95.000 95.535 98.530 ;
        RECT 95.970 98.525 96.285 98.530 ;
        RECT 95.970 95.000 96.200 98.525 ;
        RECT 95.340 94.565 96.200 95.000 ;
        RECT 91.200 94.340 92.290 94.550 ;
        RECT 91.200 94.240 92.160 94.340 ;
        RECT 93.080 94.335 94.040 94.565 ;
        RECT 94.960 94.340 96.200 94.565 ;
        RECT 94.960 94.335 95.920 94.340 ;
        RECT 96.700 93.770 97.890 95.930 ;
        RECT 98.360 93.770 99.550 95.930 ;
        RECT 101.540 94.960 101.890 97.180 ;
        RECT 107.940 94.770 108.170 98.530 ;
        RECT 108.605 94.565 108.795 98.975 ;
        RECT 109.385 98.770 109.925 99.270 ;
        RECT 110.110 99.205 111.050 99.515 ;
        RECT 110.100 98.975 111.060 99.205 ;
        RECT 109.230 98.535 110.050 98.770 ;
        RECT 109.230 98.530 109.575 98.535 ;
        RECT 109.230 95.010 109.460 98.530 ;
        RECT 109.820 95.010 110.050 98.535 ;
        RECT 109.230 94.820 110.050 95.010 ;
        RECT 109.230 94.770 109.460 94.820 ;
        RECT 109.820 94.770 110.050 94.820 ;
        RECT 110.485 94.565 110.675 98.975 ;
        RECT 111.235 98.770 111.425 99.950 ;
        RECT 111.110 98.525 111.425 98.770 ;
        RECT 111.595 99.950 111.930 100.185 ;
        RECT 111.595 98.770 111.785 99.950 ;
        RECT 112.365 99.750 112.555 104.155 ;
        RECT 114.240 103.720 115.195 104.155 ;
        RECT 114.245 100.190 114.435 103.720 ;
        RECT 114.870 103.710 115.195 103.720 ;
        RECT 114.870 100.190 115.100 103.710 ;
        RECT 114.245 100.185 115.180 100.190 ;
        RECT 114.245 100.180 115.185 100.185 ;
        RECT 114.240 99.750 115.185 100.180 ;
        RECT 116.125 99.750 116.315 104.155 ;
        RECT 118.000 104.010 118.830 104.155 ;
        RECT 116.560 103.410 117.170 104.010 ;
        RECT 118.000 103.720 119.050 104.010 ;
        RECT 116.750 100.155 116.980 103.410 ;
        RECT 118.005 100.190 118.195 103.720 ;
        RECT 118.440 103.410 119.050 103.720 ;
        RECT 118.630 100.195 118.860 103.410 ;
        RECT 119.420 102.045 119.670 104.710 ;
        RECT 120.190 102.020 121.380 104.180 ;
        RECT 124.200 102.750 124.550 104.970 ;
        RECT 118.630 100.190 118.945 100.195 ;
        RECT 116.750 99.950 117.065 100.155 ;
        RECT 111.980 98.970 112.940 99.750 ;
        RECT 113.860 98.970 115.185 99.750 ;
        RECT 115.720 98.970 116.720 99.750 ;
        RECT 111.595 98.530 111.930 98.770 ;
        RECT 111.110 94.770 111.340 98.525 ;
        RECT 111.700 94.770 111.930 98.530 ;
        RECT 112.365 94.570 112.555 98.970 ;
        RECT 114.245 98.525 115.185 98.970 ;
        RECT 114.245 98.520 115.180 98.525 ;
        RECT 114.245 95.000 114.435 98.520 ;
        RECT 114.870 95.000 115.100 98.520 ;
        RECT 114.245 94.770 115.100 95.000 ;
        RECT 114.245 94.570 115.070 94.770 ;
        RECT 108.220 94.335 109.180 94.565 ;
        RECT 110.100 94.335 111.060 94.565 ;
        RECT 111.980 94.240 112.940 94.570 ;
        RECT 113.860 94.550 115.070 94.570 ;
        RECT 116.125 94.565 116.315 98.970 ;
        RECT 116.875 98.770 117.065 99.950 ;
        RECT 118.005 99.750 118.945 100.190 ;
        RECT 117.600 98.970 118.945 99.750 ;
        RECT 124.200 99.460 124.550 101.680 ;
        RECT 116.750 98.530 117.065 98.770 ;
        RECT 118.005 98.530 118.945 98.970 ;
        RECT 116.750 94.770 116.980 98.530 ;
        RECT 118.005 95.000 118.195 98.530 ;
        RECT 118.630 98.525 118.945 98.530 ;
        RECT 118.630 95.000 118.860 98.525 ;
        RECT 118.000 94.565 118.860 95.000 ;
        RECT 113.860 94.340 114.950 94.550 ;
        RECT 113.860 94.240 114.820 94.340 ;
        RECT 115.740 94.335 116.700 94.565 ;
        RECT 117.620 94.340 118.860 94.565 ;
        RECT 117.620 94.335 118.580 94.340 ;
        RECT 119.360 93.770 120.550 95.930 ;
        RECT 121.020 93.770 122.210 95.930 ;
        RECT 124.200 94.960 124.550 97.180 ;
        RECT 40.270 93.240 41.170 93.290 ;
        RECT 42.150 93.240 43.050 93.290 ;
        RECT 40.240 93.010 41.200 93.240 ;
        RECT 42.120 93.215 43.080 93.240 ;
        RECT 42.120 93.010 43.340 93.215 ;
        RECT 44.000 93.010 44.960 93.240 ;
        RECT 45.880 93.010 46.840 93.240 ;
        RECT 47.740 93.010 48.740 93.330 ;
        RECT 49.620 93.010 50.620 93.330 ;
        RECT 51.500 93.240 52.500 93.330 ;
        RECT 62.930 93.240 63.830 93.290 ;
        RECT 64.810 93.240 65.710 93.290 ;
        RECT 51.500 93.010 52.760 93.240 ;
        RECT 62.900 93.010 63.860 93.240 ;
        RECT 64.780 93.215 65.740 93.240 ;
        RECT 64.780 93.010 66.000 93.215 ;
        RECT 66.660 93.010 67.620 93.240 ;
        RECT 68.540 93.010 69.500 93.240 ;
        RECT 70.400 93.010 71.400 93.330 ;
        RECT 72.280 93.010 73.280 93.330 ;
        RECT 74.160 93.240 75.160 93.330 ;
        RECT 85.590 93.240 86.490 93.290 ;
        RECT 87.470 93.240 88.370 93.290 ;
        RECT 74.160 93.010 75.420 93.240 ;
        RECT 85.560 93.010 86.520 93.240 ;
        RECT 87.440 93.215 88.400 93.240 ;
        RECT 87.440 93.010 88.660 93.215 ;
        RECT 89.320 93.010 90.280 93.240 ;
        RECT 91.200 93.010 92.160 93.240 ;
        RECT 93.060 93.010 94.060 93.330 ;
        RECT 94.940 93.010 95.940 93.330 ;
        RECT 96.820 93.240 97.820 93.330 ;
        RECT 108.250 93.240 109.150 93.290 ;
        RECT 110.130 93.240 111.030 93.290 ;
        RECT 96.820 93.010 98.080 93.240 ;
        RECT 108.220 93.010 109.180 93.240 ;
        RECT 110.100 93.215 111.060 93.240 ;
        RECT 110.100 93.010 111.320 93.215 ;
        RECT 111.980 93.010 112.940 93.240 ;
        RECT 113.860 93.010 114.820 93.240 ;
        RECT 115.720 93.010 116.720 93.330 ;
        RECT 117.600 93.010 118.600 93.330 ;
        RECT 119.480 93.240 120.480 93.330 ;
        RECT 119.480 93.010 120.740 93.240 ;
        RECT 40.270 92.970 41.170 93.010 ;
        RECT 42.150 92.970 43.340 93.010 ;
        RECT 39.960 91.085 40.190 92.850 ;
        RECT 39.875 90.850 40.190 91.085 ;
        RECT 39.875 89.760 40.065 90.850 ;
        RECT 40.625 90.690 40.815 92.970 ;
        RECT 42.500 92.850 43.340 92.970 ;
        RECT 42.500 92.620 43.360 92.850 ;
        RECT 42.505 91.090 42.695 92.620 ;
        RECT 43.130 91.095 43.360 92.620 ;
        RECT 43.720 91.105 43.950 92.850 ;
        RECT 43.130 91.090 43.455 91.095 ;
        RECT 42.505 90.690 43.455 91.090 ;
        RECT 40.240 89.920 41.200 90.690 ;
        RECT 36.200 89.135 36.530 89.540 ;
        RECT 36.800 89.135 37.130 89.540 ;
        RECT 37.400 89.135 37.730 89.540 ;
        RECT 38.000 89.135 38.330 89.540 ;
        RECT 39.875 89.520 40.190 89.760 ;
        RECT 34.875 88.885 38.330 89.135 ;
        RECT 34.875 86.600 35.125 88.885 ;
        RECT 36.200 88.480 36.530 88.885 ;
        RECT 36.800 88.480 37.130 88.885 ;
        RECT 37.400 88.480 37.730 88.885 ;
        RECT 38.000 88.480 38.330 88.885 ;
        RECT 39.960 88.370 40.190 89.520 ;
        RECT 36.270 87.620 36.730 87.850 ;
        RECT 37.670 87.620 38.130 87.850 ;
        RECT 39.820 87.760 40.420 88.370 ;
        RECT 35.990 87.115 36.220 87.460 ;
        RECT 35.825 86.960 36.220 87.115 ;
        RECT 35.825 86.925 36.205 86.960 ;
        RECT 35.825 86.600 36.015 86.925 ;
        RECT 36.405 86.800 36.595 87.620 ;
        RECT 37.390 87.115 37.620 87.460 ;
        RECT 37.225 86.960 37.620 87.115 ;
        RECT 37.225 86.925 37.605 86.960 ;
        RECT 34.840 85.825 36.015 86.600 ;
        RECT 36.270 86.730 36.730 86.800 ;
        RECT 36.270 86.570 36.755 86.730 ;
        RECT 36.405 86.505 36.755 86.570 ;
        RECT 37.225 86.505 37.415 86.925 ;
        RECT 37.805 86.800 37.995 87.620 ;
        RECT 37.670 86.670 38.130 86.800 ;
        RECT 37.670 86.570 38.150 86.670 ;
        RECT 39.820 86.610 40.015 87.760 ;
        RECT 40.625 87.600 40.815 89.920 ;
        RECT 42.120 89.910 43.455 90.690 ;
        RECT 42.505 89.520 43.455 89.910 ;
        RECT 43.635 90.850 43.950 91.105 ;
        RECT 43.635 89.760 43.825 90.850 ;
        RECT 44.385 90.690 44.575 93.010 ;
        RECT 45.010 92.800 45.240 92.850 ;
        RECT 45.600 92.800 45.830 92.850 ;
        RECT 45.010 92.610 45.830 92.800 ;
        RECT 45.010 91.090 45.240 92.610 ;
        RECT 45.600 91.090 45.830 92.610 ;
        RECT 45.010 90.850 45.830 91.090 ;
        RECT 44.000 89.920 44.960 90.690 ;
        RECT 43.635 89.520 43.950 89.760 ;
        RECT 42.505 88.010 42.695 89.520 ;
        RECT 43.130 88.010 43.360 89.520 ;
        RECT 43.720 88.370 43.950 89.520 ;
        RECT 42.500 88.005 43.440 88.010 ;
        RECT 42.500 87.600 43.445 88.005 ;
        RECT 40.240 87.580 41.200 87.600 ;
        RECT 42.120 87.580 43.445 87.600 ;
        RECT 40.240 87.390 43.445 87.580 ;
        RECT 40.240 87.370 41.200 87.390 ;
        RECT 42.120 87.370 43.445 87.390 ;
        RECT 40.240 86.815 41.200 87.045 ;
        RECT 42.120 86.815 43.080 87.045 ;
        RECT 36.405 86.315 37.415 86.505 ;
        RECT 36.405 86.235 36.755 86.315 ;
        RECT 36.270 86.155 36.755 86.235 ;
        RECT 36.270 86.005 36.730 86.155 ;
        RECT 34.840 85.800 36.200 85.825 ;
        RECT 34.840 85.600 36.220 85.800 ;
        RECT 35.990 84.800 36.220 85.600 ;
        RECT 36.405 84.595 36.595 86.005 ;
        RECT 37.225 85.825 37.415 86.315 ;
        RECT 37.805 86.515 38.150 86.570 ;
        RECT 38.590 86.515 39.590 86.600 ;
        RECT 37.805 86.325 39.590 86.515 ;
        RECT 37.805 86.235 38.150 86.325 ;
        RECT 37.670 86.200 38.150 86.235 ;
        RECT 37.670 86.005 38.130 86.200 ;
        RECT 37.225 85.800 37.605 85.825 ;
        RECT 37.225 85.635 37.620 85.800 ;
        RECT 37.390 84.800 37.620 85.635 ;
        RECT 37.805 84.595 37.995 86.005 ;
        RECT 38.590 85.600 39.590 86.325 ;
        RECT 39.820 86.010 40.420 86.610 ;
        RECT 36.270 84.365 36.730 84.595 ;
        RECT 37.670 84.365 38.130 84.595 ;
        RECT 39.960 82.855 40.190 86.010 ;
        RECT 39.875 82.610 40.190 82.855 ;
        RECT 39.875 81.430 40.065 82.610 ;
        RECT 40.625 82.405 40.815 86.815 ;
        RECT 41.250 86.560 41.480 86.610 ;
        RECT 41.840 86.560 42.070 86.610 ;
        RECT 41.250 86.370 42.070 86.560 ;
        RECT 41.250 82.855 41.480 86.370 ;
        RECT 41.250 82.850 41.595 82.855 ;
        RECT 41.840 82.850 42.070 86.370 ;
        RECT 41.250 82.610 42.070 82.850 ;
        RECT 40.240 82.175 41.200 82.405 ;
        RECT 40.300 81.865 41.140 82.175 ;
        RECT 41.405 82.120 41.945 82.610 ;
        RECT 42.505 82.405 42.695 86.815 ;
        RECT 43.255 86.610 43.445 87.370 ;
        RECT 43.130 86.365 43.445 86.610 ;
        RECT 43.620 87.770 44.230 88.370 ;
        RECT 43.620 87.760 43.950 87.770 ;
        RECT 43.620 86.610 43.810 87.760 ;
        RECT 44.385 87.600 44.575 89.920 ;
        RECT 45.145 89.760 45.705 90.850 ;
        RECT 46.265 90.690 46.455 93.010 ;
        RECT 46.890 91.090 47.120 92.850 ;
        RECT 46.890 90.850 47.205 91.090 ;
        RECT 45.880 89.920 46.840 90.690 ;
        RECT 45.010 89.520 45.830 89.760 ;
        RECT 45.010 88.000 45.240 89.520 ;
        RECT 45.600 88.000 45.830 89.520 ;
        RECT 45.010 87.810 45.830 88.000 ;
        RECT 45.010 87.760 45.240 87.810 ;
        RECT 45.600 87.760 45.830 87.810 ;
        RECT 46.265 87.600 46.455 89.920 ;
        RECT 47.015 89.760 47.205 90.850 ;
        RECT 48.145 90.690 48.335 93.010 ;
        RECT 48.770 91.095 49.000 92.850 ;
        RECT 48.770 90.850 49.085 91.095 ;
        RECT 47.740 89.920 48.740 90.690 ;
        RECT 46.890 89.515 47.205 89.760 ;
        RECT 46.890 88.005 47.120 89.515 ;
        RECT 46.890 87.760 47.215 88.005 ;
        RECT 44.000 87.370 44.960 87.600 ;
        RECT 45.880 87.370 46.840 87.600 ;
        RECT 47.025 87.050 47.215 87.760 ;
        RECT 48.145 87.600 48.335 89.920 ;
        RECT 48.895 89.760 49.085 90.850 ;
        RECT 50.025 90.690 50.215 93.010 ;
        RECT 50.650 91.105 50.880 92.850 ;
        RECT 51.900 92.610 52.760 93.010 ;
        RECT 62.930 92.970 63.830 93.010 ;
        RECT 64.810 92.970 66.000 93.010 ;
        RECT 50.650 90.850 50.965 91.105 ;
        RECT 49.620 89.920 50.620 90.690 ;
        RECT 48.770 89.515 49.085 89.760 ;
        RECT 48.770 88.370 49.000 89.515 ;
        RECT 48.590 87.770 49.190 88.370 ;
        RECT 48.770 87.760 49.000 87.770 ;
        RECT 50.025 87.600 50.215 89.920 ;
        RECT 50.775 89.760 50.965 90.850 ;
        RECT 51.900 91.080 52.095 92.610 ;
        RECT 52.530 91.090 52.760 92.610 ;
        RECT 52.530 91.080 52.855 91.090 ;
        RECT 51.900 90.690 52.855 91.080 ;
        RECT 51.500 89.920 52.855 90.690 ;
        RECT 53.410 90.355 54.060 90.540 ;
        RECT 55.010 90.355 55.330 90.390 ;
        RECT 53.410 90.165 55.330 90.355 ;
        RECT 53.410 89.990 54.060 90.165 ;
        RECT 55.010 90.130 55.330 90.165 ;
        RECT 50.650 89.520 50.965 89.760 ;
        RECT 50.650 88.370 50.880 89.520 ;
        RECT 51.900 89.515 52.855 89.920 ;
        RECT 56.220 89.910 56.570 92.130 ;
        RECT 62.620 91.085 62.850 92.850 ;
        RECT 62.535 90.850 62.850 91.085 ;
        RECT 62.535 89.760 62.725 90.850 ;
        RECT 63.285 90.690 63.475 92.970 ;
        RECT 65.160 92.850 66.000 92.970 ;
        RECT 65.160 92.620 66.020 92.850 ;
        RECT 65.165 91.090 65.355 92.620 ;
        RECT 65.790 91.095 66.020 92.620 ;
        RECT 66.380 91.105 66.610 92.850 ;
        RECT 65.790 91.090 66.115 91.095 ;
        RECT 65.165 90.690 66.115 91.090 ;
        RECT 62.900 89.920 63.860 90.690 ;
        RECT 51.900 89.510 52.850 89.515 ;
        RECT 50.470 87.770 51.070 88.370 ;
        RECT 51.900 87.990 52.095 89.510 ;
        RECT 52.530 87.990 52.760 89.510 ;
        RECT 58.860 89.135 59.190 89.540 ;
        RECT 59.460 89.135 59.790 89.540 ;
        RECT 60.060 89.135 60.390 89.540 ;
        RECT 60.660 89.135 60.990 89.540 ;
        RECT 62.535 89.520 62.850 89.760 ;
        RECT 50.650 87.760 50.880 87.770 ;
        RECT 51.900 87.600 52.760 87.990 ;
        RECT 57.535 88.885 60.990 89.135 ;
        RECT 47.740 87.370 52.760 87.600 ;
        RECT 44.000 86.820 47.215 87.050 ;
        RECT 44.000 86.815 44.960 86.820 ;
        RECT 45.880 86.815 47.215 86.820 ;
        RECT 47.760 86.815 48.720 87.045 ;
        RECT 49.640 87.010 50.600 87.045 ;
        RECT 49.640 86.815 50.850 87.010 ;
        RECT 43.620 86.600 43.950 86.610 ;
        RECT 43.130 82.845 43.360 86.365 ;
        RECT 43.620 86.000 44.230 86.600 ;
        RECT 43.720 82.845 43.950 86.000 ;
        RECT 43.130 82.610 43.445 82.845 ;
        RECT 42.120 82.175 43.080 82.405 ;
        RECT 41.395 81.930 41.945 82.120 ;
        RECT 40.240 81.635 41.200 81.865 ;
        RECT 39.875 81.190 40.190 81.430 ;
        RECT 39.960 77.430 40.190 81.190 ;
        RECT 40.625 77.225 40.815 81.635 ;
        RECT 41.405 81.430 41.945 81.930 ;
        RECT 42.130 81.865 43.070 82.175 ;
        RECT 42.120 81.635 43.080 81.865 ;
        RECT 41.250 81.195 42.070 81.430 ;
        RECT 41.250 81.190 41.595 81.195 ;
        RECT 41.250 77.670 41.480 81.190 ;
        RECT 41.840 77.670 42.070 81.195 ;
        RECT 41.250 77.480 42.070 77.670 ;
        RECT 41.250 77.430 41.480 77.480 ;
        RECT 41.840 77.430 42.070 77.480 ;
        RECT 42.505 77.225 42.695 81.635 ;
        RECT 43.255 81.430 43.445 82.610 ;
        RECT 43.130 81.185 43.445 81.430 ;
        RECT 43.615 82.610 43.950 82.845 ;
        RECT 43.615 81.430 43.805 82.610 ;
        RECT 44.385 82.410 44.575 86.815 ;
        RECT 46.260 86.380 47.215 86.815 ;
        RECT 46.265 82.850 46.455 86.380 ;
        RECT 46.890 86.370 47.215 86.380 ;
        RECT 46.890 82.850 47.120 86.370 ;
        RECT 46.265 82.845 47.200 82.850 ;
        RECT 46.265 82.840 47.205 82.845 ;
        RECT 46.260 82.410 47.205 82.840 ;
        RECT 48.145 82.410 48.335 86.815 ;
        RECT 50.020 86.670 50.850 86.815 ;
        RECT 48.580 86.070 49.190 86.670 ;
        RECT 50.020 86.380 51.070 86.670 ;
        RECT 48.770 82.815 49.000 86.070 ;
        RECT 50.025 82.850 50.215 86.380 ;
        RECT 50.460 86.070 51.070 86.380 ;
        RECT 50.650 82.855 50.880 86.070 ;
        RECT 51.440 84.705 51.690 87.370 ;
        RECT 52.210 84.680 53.400 86.840 ;
        RECT 56.220 85.410 56.570 87.630 ;
        RECT 57.535 86.600 57.785 88.885 ;
        RECT 58.860 88.480 59.190 88.885 ;
        RECT 59.460 88.480 59.790 88.885 ;
        RECT 60.060 88.480 60.390 88.885 ;
        RECT 60.660 88.480 60.990 88.885 ;
        RECT 62.620 88.370 62.850 89.520 ;
        RECT 58.930 87.620 59.390 87.850 ;
        RECT 60.330 87.620 60.790 87.850 ;
        RECT 62.480 87.760 63.080 88.370 ;
        RECT 58.650 87.115 58.880 87.460 ;
        RECT 58.485 86.960 58.880 87.115 ;
        RECT 58.485 86.925 58.865 86.960 ;
        RECT 58.485 86.600 58.675 86.925 ;
        RECT 59.065 86.800 59.255 87.620 ;
        RECT 60.050 87.115 60.280 87.460 ;
        RECT 59.885 86.960 60.280 87.115 ;
        RECT 59.885 86.925 60.265 86.960 ;
        RECT 57.500 85.825 58.675 86.600 ;
        RECT 58.930 86.730 59.390 86.800 ;
        RECT 58.930 86.570 59.415 86.730 ;
        RECT 59.065 86.505 59.415 86.570 ;
        RECT 59.885 86.505 60.075 86.925 ;
        RECT 60.465 86.800 60.655 87.620 ;
        RECT 60.330 86.670 60.790 86.800 ;
        RECT 60.330 86.570 60.810 86.670 ;
        RECT 62.480 86.610 62.675 87.760 ;
        RECT 63.285 87.600 63.475 89.920 ;
        RECT 64.780 89.910 66.115 90.690 ;
        RECT 65.165 89.520 66.115 89.910 ;
        RECT 66.295 90.850 66.610 91.105 ;
        RECT 66.295 89.760 66.485 90.850 ;
        RECT 67.045 90.690 67.235 93.010 ;
        RECT 67.670 92.800 67.900 92.850 ;
        RECT 68.260 92.800 68.490 92.850 ;
        RECT 67.670 92.610 68.490 92.800 ;
        RECT 67.670 91.090 67.900 92.610 ;
        RECT 68.260 91.090 68.490 92.610 ;
        RECT 67.670 90.850 68.490 91.090 ;
        RECT 66.660 89.920 67.620 90.690 ;
        RECT 66.295 89.520 66.610 89.760 ;
        RECT 65.165 88.010 65.355 89.520 ;
        RECT 65.790 88.010 66.020 89.520 ;
        RECT 66.380 88.370 66.610 89.520 ;
        RECT 65.160 88.005 66.100 88.010 ;
        RECT 65.160 87.600 66.105 88.005 ;
        RECT 62.900 87.580 63.860 87.600 ;
        RECT 64.780 87.580 66.105 87.600 ;
        RECT 62.900 87.390 66.105 87.580 ;
        RECT 62.900 87.370 63.860 87.390 ;
        RECT 64.780 87.370 66.105 87.390 ;
        RECT 62.900 86.815 63.860 87.045 ;
        RECT 64.780 86.815 65.740 87.045 ;
        RECT 59.065 86.315 60.075 86.505 ;
        RECT 59.065 86.235 59.415 86.315 ;
        RECT 58.930 86.155 59.415 86.235 ;
        RECT 58.930 86.005 59.390 86.155 ;
        RECT 57.500 85.800 58.860 85.825 ;
        RECT 57.500 85.600 58.880 85.800 ;
        RECT 58.650 84.800 58.880 85.600 ;
        RECT 59.065 84.595 59.255 86.005 ;
        RECT 59.885 85.825 60.075 86.315 ;
        RECT 60.465 86.515 60.810 86.570 ;
        RECT 61.250 86.515 62.250 86.600 ;
        RECT 60.465 86.325 62.250 86.515 ;
        RECT 60.465 86.235 60.810 86.325 ;
        RECT 60.330 86.200 60.810 86.235 ;
        RECT 60.330 86.005 60.790 86.200 ;
        RECT 59.885 85.800 60.265 85.825 ;
        RECT 59.885 85.635 60.280 85.800 ;
        RECT 60.050 84.800 60.280 85.635 ;
        RECT 60.465 84.595 60.655 86.005 ;
        RECT 61.250 85.600 62.250 86.325 ;
        RECT 62.480 86.010 63.080 86.610 ;
        RECT 58.930 84.365 59.390 84.595 ;
        RECT 60.330 84.365 60.790 84.595 ;
        RECT 50.650 82.850 50.965 82.855 ;
        RECT 48.770 82.610 49.085 82.815 ;
        RECT 44.000 81.630 44.960 82.410 ;
        RECT 45.880 81.630 47.205 82.410 ;
        RECT 47.740 81.630 48.740 82.410 ;
        RECT 43.615 81.190 43.950 81.430 ;
        RECT 43.130 77.430 43.360 81.185 ;
        RECT 43.720 77.430 43.950 81.190 ;
        RECT 44.385 77.230 44.575 81.630 ;
        RECT 46.265 81.185 47.205 81.630 ;
        RECT 46.265 81.180 47.200 81.185 ;
        RECT 46.265 77.660 46.455 81.180 ;
        RECT 46.890 77.660 47.120 81.180 ;
        RECT 46.265 77.430 47.120 77.660 ;
        RECT 46.265 77.230 47.090 77.430 ;
        RECT 40.240 76.995 41.200 77.225 ;
        RECT 42.120 76.995 43.080 77.225 ;
        RECT 44.000 76.900 44.960 77.230 ;
        RECT 45.880 77.210 47.090 77.230 ;
        RECT 48.145 77.225 48.335 81.630 ;
        RECT 48.895 81.430 49.085 82.610 ;
        RECT 50.025 82.410 50.965 82.850 ;
        RECT 49.620 81.630 50.965 82.410 ;
        RECT 56.220 82.120 56.570 84.340 ;
        RECT 62.620 82.855 62.850 86.010 ;
        RECT 62.535 82.610 62.850 82.855 ;
        RECT 48.770 81.190 49.085 81.430 ;
        RECT 50.025 81.190 50.965 81.630 ;
        RECT 62.535 81.430 62.725 82.610 ;
        RECT 63.285 82.405 63.475 86.815 ;
        RECT 63.910 86.560 64.140 86.610 ;
        RECT 64.500 86.560 64.730 86.610 ;
        RECT 63.910 86.370 64.730 86.560 ;
        RECT 63.910 82.855 64.140 86.370 ;
        RECT 63.910 82.850 64.255 82.855 ;
        RECT 64.500 82.850 64.730 86.370 ;
        RECT 63.910 82.610 64.730 82.850 ;
        RECT 62.900 82.175 63.860 82.405 ;
        RECT 62.960 81.865 63.800 82.175 ;
        RECT 64.065 82.120 64.605 82.610 ;
        RECT 65.165 82.405 65.355 86.815 ;
        RECT 65.915 86.610 66.105 87.370 ;
        RECT 65.790 86.365 66.105 86.610 ;
        RECT 66.280 87.770 66.890 88.370 ;
        RECT 66.280 87.760 66.610 87.770 ;
        RECT 66.280 86.610 66.470 87.760 ;
        RECT 67.045 87.600 67.235 89.920 ;
        RECT 67.805 89.760 68.365 90.850 ;
        RECT 68.925 90.690 69.115 93.010 ;
        RECT 69.550 91.090 69.780 92.850 ;
        RECT 69.550 90.850 69.865 91.090 ;
        RECT 68.540 89.920 69.500 90.690 ;
        RECT 67.670 89.520 68.490 89.760 ;
        RECT 67.670 88.000 67.900 89.520 ;
        RECT 68.260 88.000 68.490 89.520 ;
        RECT 67.670 87.810 68.490 88.000 ;
        RECT 67.670 87.760 67.900 87.810 ;
        RECT 68.260 87.760 68.490 87.810 ;
        RECT 68.925 87.600 69.115 89.920 ;
        RECT 69.675 89.760 69.865 90.850 ;
        RECT 70.805 90.690 70.995 93.010 ;
        RECT 71.430 91.095 71.660 92.850 ;
        RECT 71.430 90.850 71.745 91.095 ;
        RECT 70.400 89.920 71.400 90.690 ;
        RECT 69.550 89.515 69.865 89.760 ;
        RECT 69.550 88.005 69.780 89.515 ;
        RECT 69.550 87.760 69.875 88.005 ;
        RECT 66.660 87.370 67.620 87.600 ;
        RECT 68.540 87.370 69.500 87.600 ;
        RECT 69.685 87.050 69.875 87.760 ;
        RECT 70.805 87.600 70.995 89.920 ;
        RECT 71.555 89.760 71.745 90.850 ;
        RECT 72.685 90.690 72.875 93.010 ;
        RECT 73.310 91.105 73.540 92.850 ;
        RECT 74.560 92.610 75.420 93.010 ;
        RECT 85.590 92.970 86.490 93.010 ;
        RECT 87.470 92.970 88.660 93.010 ;
        RECT 73.310 90.850 73.625 91.105 ;
        RECT 72.280 89.920 73.280 90.690 ;
        RECT 71.430 89.515 71.745 89.760 ;
        RECT 71.430 88.370 71.660 89.515 ;
        RECT 71.250 87.770 71.850 88.370 ;
        RECT 71.430 87.760 71.660 87.770 ;
        RECT 72.685 87.600 72.875 89.920 ;
        RECT 73.435 89.760 73.625 90.850 ;
        RECT 74.560 91.080 74.755 92.610 ;
        RECT 75.190 91.090 75.420 92.610 ;
        RECT 75.190 91.080 75.515 91.090 ;
        RECT 74.560 90.690 75.515 91.080 ;
        RECT 74.160 89.920 75.515 90.690 ;
        RECT 76.070 90.355 76.720 90.540 ;
        RECT 77.670 90.355 77.990 90.390 ;
        RECT 76.070 90.165 77.990 90.355 ;
        RECT 76.070 89.990 76.720 90.165 ;
        RECT 77.670 90.130 77.990 90.165 ;
        RECT 73.310 89.520 73.625 89.760 ;
        RECT 73.310 88.370 73.540 89.520 ;
        RECT 74.560 89.515 75.515 89.920 ;
        RECT 78.880 89.910 79.230 92.130 ;
        RECT 85.280 91.085 85.510 92.850 ;
        RECT 85.195 90.850 85.510 91.085 ;
        RECT 85.195 89.760 85.385 90.850 ;
        RECT 85.945 90.690 86.135 92.970 ;
        RECT 87.820 92.850 88.660 92.970 ;
        RECT 87.820 92.620 88.680 92.850 ;
        RECT 87.825 91.090 88.015 92.620 ;
        RECT 88.450 91.095 88.680 92.620 ;
        RECT 89.040 91.105 89.270 92.850 ;
        RECT 88.450 91.090 88.775 91.095 ;
        RECT 87.825 90.690 88.775 91.090 ;
        RECT 85.560 89.920 86.520 90.690 ;
        RECT 74.560 89.510 75.510 89.515 ;
        RECT 73.130 87.770 73.730 88.370 ;
        RECT 74.560 87.990 74.755 89.510 ;
        RECT 75.190 87.990 75.420 89.510 ;
        RECT 81.520 89.135 81.850 89.540 ;
        RECT 82.120 89.135 82.450 89.540 ;
        RECT 82.720 89.135 83.050 89.540 ;
        RECT 83.320 89.135 83.650 89.540 ;
        RECT 85.195 89.520 85.510 89.760 ;
        RECT 73.310 87.760 73.540 87.770 ;
        RECT 74.560 87.600 75.420 87.990 ;
        RECT 80.195 88.885 83.650 89.135 ;
        RECT 70.400 87.370 75.420 87.600 ;
        RECT 66.660 86.820 69.875 87.050 ;
        RECT 66.660 86.815 67.620 86.820 ;
        RECT 68.540 86.815 69.875 86.820 ;
        RECT 70.420 86.815 71.380 87.045 ;
        RECT 72.300 87.010 73.260 87.045 ;
        RECT 72.300 86.815 73.510 87.010 ;
        RECT 66.280 86.600 66.610 86.610 ;
        RECT 65.790 82.845 66.020 86.365 ;
        RECT 66.280 86.000 66.890 86.600 ;
        RECT 66.380 82.845 66.610 86.000 ;
        RECT 65.790 82.610 66.105 82.845 ;
        RECT 64.780 82.175 65.740 82.405 ;
        RECT 64.055 81.930 64.605 82.120 ;
        RECT 62.900 81.635 63.860 81.865 ;
        RECT 62.535 81.190 62.850 81.430 ;
        RECT 48.770 77.430 49.000 81.190 ;
        RECT 50.025 77.660 50.215 81.190 ;
        RECT 50.650 81.185 50.965 81.190 ;
        RECT 50.650 77.660 50.880 81.185 ;
        RECT 50.020 77.225 50.880 77.660 ;
        RECT 45.880 77.000 46.970 77.210 ;
        RECT 45.880 76.900 46.840 77.000 ;
        RECT 47.760 76.995 48.720 77.225 ;
        RECT 49.640 77.000 50.880 77.225 ;
        RECT 49.640 76.995 50.600 77.000 ;
        RECT 51.380 76.430 52.570 78.590 ;
        RECT 53.040 76.430 54.230 78.590 ;
        RECT 56.220 77.620 56.570 79.840 ;
        RECT 62.620 77.430 62.850 81.190 ;
        RECT 63.285 77.225 63.475 81.635 ;
        RECT 64.065 81.430 64.605 81.930 ;
        RECT 64.790 81.865 65.730 82.175 ;
        RECT 64.780 81.635 65.740 81.865 ;
        RECT 63.910 81.195 64.730 81.430 ;
        RECT 63.910 81.190 64.255 81.195 ;
        RECT 63.910 77.670 64.140 81.190 ;
        RECT 64.500 77.670 64.730 81.195 ;
        RECT 63.910 77.480 64.730 77.670 ;
        RECT 63.910 77.430 64.140 77.480 ;
        RECT 64.500 77.430 64.730 77.480 ;
        RECT 65.165 77.225 65.355 81.635 ;
        RECT 65.915 81.430 66.105 82.610 ;
        RECT 65.790 81.185 66.105 81.430 ;
        RECT 66.275 82.610 66.610 82.845 ;
        RECT 66.275 81.430 66.465 82.610 ;
        RECT 67.045 82.410 67.235 86.815 ;
        RECT 68.920 86.380 69.875 86.815 ;
        RECT 68.925 82.850 69.115 86.380 ;
        RECT 69.550 86.370 69.875 86.380 ;
        RECT 69.550 82.850 69.780 86.370 ;
        RECT 68.925 82.845 69.860 82.850 ;
        RECT 68.925 82.840 69.865 82.845 ;
        RECT 68.920 82.410 69.865 82.840 ;
        RECT 70.805 82.410 70.995 86.815 ;
        RECT 72.680 86.670 73.510 86.815 ;
        RECT 71.240 86.070 71.850 86.670 ;
        RECT 72.680 86.380 73.730 86.670 ;
        RECT 71.430 82.815 71.660 86.070 ;
        RECT 72.685 82.850 72.875 86.380 ;
        RECT 73.120 86.070 73.730 86.380 ;
        RECT 73.310 82.855 73.540 86.070 ;
        RECT 74.100 84.705 74.350 87.370 ;
        RECT 74.870 84.680 76.060 86.840 ;
        RECT 78.880 85.410 79.230 87.630 ;
        RECT 80.195 86.600 80.445 88.885 ;
        RECT 81.520 88.480 81.850 88.885 ;
        RECT 82.120 88.480 82.450 88.885 ;
        RECT 82.720 88.480 83.050 88.885 ;
        RECT 83.320 88.480 83.650 88.885 ;
        RECT 85.280 88.370 85.510 89.520 ;
        RECT 81.590 87.620 82.050 87.850 ;
        RECT 82.990 87.620 83.450 87.850 ;
        RECT 85.140 87.760 85.740 88.370 ;
        RECT 81.310 87.115 81.540 87.460 ;
        RECT 81.145 86.960 81.540 87.115 ;
        RECT 81.145 86.925 81.525 86.960 ;
        RECT 81.145 86.600 81.335 86.925 ;
        RECT 81.725 86.800 81.915 87.620 ;
        RECT 82.710 87.115 82.940 87.460 ;
        RECT 82.545 86.960 82.940 87.115 ;
        RECT 82.545 86.925 82.925 86.960 ;
        RECT 80.160 85.825 81.335 86.600 ;
        RECT 81.590 86.730 82.050 86.800 ;
        RECT 81.590 86.570 82.075 86.730 ;
        RECT 81.725 86.505 82.075 86.570 ;
        RECT 82.545 86.505 82.735 86.925 ;
        RECT 83.125 86.800 83.315 87.620 ;
        RECT 82.990 86.670 83.450 86.800 ;
        RECT 82.990 86.570 83.470 86.670 ;
        RECT 85.140 86.610 85.335 87.760 ;
        RECT 85.945 87.600 86.135 89.920 ;
        RECT 87.440 89.910 88.775 90.690 ;
        RECT 87.825 89.520 88.775 89.910 ;
        RECT 88.955 90.850 89.270 91.105 ;
        RECT 88.955 89.760 89.145 90.850 ;
        RECT 89.705 90.690 89.895 93.010 ;
        RECT 90.330 92.800 90.560 92.850 ;
        RECT 90.920 92.800 91.150 92.850 ;
        RECT 90.330 92.610 91.150 92.800 ;
        RECT 90.330 91.090 90.560 92.610 ;
        RECT 90.920 91.090 91.150 92.610 ;
        RECT 90.330 90.850 91.150 91.090 ;
        RECT 89.320 89.920 90.280 90.690 ;
        RECT 88.955 89.520 89.270 89.760 ;
        RECT 87.825 88.010 88.015 89.520 ;
        RECT 88.450 88.010 88.680 89.520 ;
        RECT 89.040 88.370 89.270 89.520 ;
        RECT 87.820 88.005 88.760 88.010 ;
        RECT 87.820 87.600 88.765 88.005 ;
        RECT 85.560 87.580 86.520 87.600 ;
        RECT 87.440 87.580 88.765 87.600 ;
        RECT 85.560 87.390 88.765 87.580 ;
        RECT 85.560 87.370 86.520 87.390 ;
        RECT 87.440 87.370 88.765 87.390 ;
        RECT 85.560 86.815 86.520 87.045 ;
        RECT 87.440 86.815 88.400 87.045 ;
        RECT 81.725 86.315 82.735 86.505 ;
        RECT 81.725 86.235 82.075 86.315 ;
        RECT 81.590 86.155 82.075 86.235 ;
        RECT 81.590 86.005 82.050 86.155 ;
        RECT 80.160 85.800 81.520 85.825 ;
        RECT 80.160 85.600 81.540 85.800 ;
        RECT 81.310 84.800 81.540 85.600 ;
        RECT 81.725 84.595 81.915 86.005 ;
        RECT 82.545 85.825 82.735 86.315 ;
        RECT 83.125 86.515 83.470 86.570 ;
        RECT 83.910 86.515 84.910 86.600 ;
        RECT 83.125 86.325 84.910 86.515 ;
        RECT 83.125 86.235 83.470 86.325 ;
        RECT 82.990 86.200 83.470 86.235 ;
        RECT 82.990 86.005 83.450 86.200 ;
        RECT 82.545 85.800 82.925 85.825 ;
        RECT 82.545 85.635 82.940 85.800 ;
        RECT 82.710 84.800 82.940 85.635 ;
        RECT 83.125 84.595 83.315 86.005 ;
        RECT 83.910 85.600 84.910 86.325 ;
        RECT 85.140 86.010 85.740 86.610 ;
        RECT 81.590 84.365 82.050 84.595 ;
        RECT 82.990 84.365 83.450 84.595 ;
        RECT 73.310 82.850 73.625 82.855 ;
        RECT 71.430 82.610 71.745 82.815 ;
        RECT 66.660 81.630 67.620 82.410 ;
        RECT 68.540 81.630 69.865 82.410 ;
        RECT 70.400 81.630 71.400 82.410 ;
        RECT 66.275 81.190 66.610 81.430 ;
        RECT 65.790 77.430 66.020 81.185 ;
        RECT 66.380 77.430 66.610 81.190 ;
        RECT 67.045 77.230 67.235 81.630 ;
        RECT 68.925 81.185 69.865 81.630 ;
        RECT 68.925 81.180 69.860 81.185 ;
        RECT 68.925 77.660 69.115 81.180 ;
        RECT 69.550 77.660 69.780 81.180 ;
        RECT 68.925 77.430 69.780 77.660 ;
        RECT 68.925 77.230 69.750 77.430 ;
        RECT 62.900 76.995 63.860 77.225 ;
        RECT 64.780 76.995 65.740 77.225 ;
        RECT 66.660 76.900 67.620 77.230 ;
        RECT 68.540 77.210 69.750 77.230 ;
        RECT 70.805 77.225 70.995 81.630 ;
        RECT 71.555 81.430 71.745 82.610 ;
        RECT 72.685 82.410 73.625 82.850 ;
        RECT 72.280 81.630 73.625 82.410 ;
        RECT 78.880 82.120 79.230 84.340 ;
        RECT 85.280 82.855 85.510 86.010 ;
        RECT 85.195 82.610 85.510 82.855 ;
        RECT 71.430 81.190 71.745 81.430 ;
        RECT 72.685 81.190 73.625 81.630 ;
        RECT 85.195 81.430 85.385 82.610 ;
        RECT 85.945 82.405 86.135 86.815 ;
        RECT 86.570 86.560 86.800 86.610 ;
        RECT 87.160 86.560 87.390 86.610 ;
        RECT 86.570 86.370 87.390 86.560 ;
        RECT 86.570 82.855 86.800 86.370 ;
        RECT 86.570 82.850 86.915 82.855 ;
        RECT 87.160 82.850 87.390 86.370 ;
        RECT 86.570 82.610 87.390 82.850 ;
        RECT 85.560 82.175 86.520 82.405 ;
        RECT 85.620 81.865 86.460 82.175 ;
        RECT 86.725 82.120 87.265 82.610 ;
        RECT 87.825 82.405 88.015 86.815 ;
        RECT 88.575 86.610 88.765 87.370 ;
        RECT 88.450 86.365 88.765 86.610 ;
        RECT 88.940 87.770 89.550 88.370 ;
        RECT 88.940 87.760 89.270 87.770 ;
        RECT 88.940 86.610 89.130 87.760 ;
        RECT 89.705 87.600 89.895 89.920 ;
        RECT 90.465 89.760 91.025 90.850 ;
        RECT 91.585 90.690 91.775 93.010 ;
        RECT 92.210 91.090 92.440 92.850 ;
        RECT 92.210 90.850 92.525 91.090 ;
        RECT 91.200 89.920 92.160 90.690 ;
        RECT 90.330 89.520 91.150 89.760 ;
        RECT 90.330 88.000 90.560 89.520 ;
        RECT 90.920 88.000 91.150 89.520 ;
        RECT 90.330 87.810 91.150 88.000 ;
        RECT 90.330 87.760 90.560 87.810 ;
        RECT 90.920 87.760 91.150 87.810 ;
        RECT 91.585 87.600 91.775 89.920 ;
        RECT 92.335 89.760 92.525 90.850 ;
        RECT 93.465 90.690 93.655 93.010 ;
        RECT 94.090 91.095 94.320 92.850 ;
        RECT 94.090 90.850 94.405 91.095 ;
        RECT 93.060 89.920 94.060 90.690 ;
        RECT 92.210 89.515 92.525 89.760 ;
        RECT 92.210 88.005 92.440 89.515 ;
        RECT 92.210 87.760 92.535 88.005 ;
        RECT 89.320 87.370 90.280 87.600 ;
        RECT 91.200 87.370 92.160 87.600 ;
        RECT 92.345 87.050 92.535 87.760 ;
        RECT 93.465 87.600 93.655 89.920 ;
        RECT 94.215 89.760 94.405 90.850 ;
        RECT 95.345 90.690 95.535 93.010 ;
        RECT 95.970 91.105 96.200 92.850 ;
        RECT 97.220 92.610 98.080 93.010 ;
        RECT 108.250 92.970 109.150 93.010 ;
        RECT 110.130 92.970 111.320 93.010 ;
        RECT 95.970 90.850 96.285 91.105 ;
        RECT 94.940 89.920 95.940 90.690 ;
        RECT 94.090 89.515 94.405 89.760 ;
        RECT 94.090 88.370 94.320 89.515 ;
        RECT 93.910 87.770 94.510 88.370 ;
        RECT 94.090 87.760 94.320 87.770 ;
        RECT 95.345 87.600 95.535 89.920 ;
        RECT 96.095 89.760 96.285 90.850 ;
        RECT 97.220 91.080 97.415 92.610 ;
        RECT 97.850 91.090 98.080 92.610 ;
        RECT 97.850 91.080 98.175 91.090 ;
        RECT 97.220 90.690 98.175 91.080 ;
        RECT 96.820 89.920 98.175 90.690 ;
        RECT 98.730 90.355 99.380 90.540 ;
        RECT 100.330 90.355 100.650 90.390 ;
        RECT 98.730 90.165 100.650 90.355 ;
        RECT 98.730 89.990 99.380 90.165 ;
        RECT 100.330 90.130 100.650 90.165 ;
        RECT 95.970 89.520 96.285 89.760 ;
        RECT 95.970 88.370 96.200 89.520 ;
        RECT 97.220 89.515 98.175 89.920 ;
        RECT 101.540 89.910 101.890 92.130 ;
        RECT 107.940 91.085 108.170 92.850 ;
        RECT 107.855 90.850 108.170 91.085 ;
        RECT 107.855 89.760 108.045 90.850 ;
        RECT 108.605 90.690 108.795 92.970 ;
        RECT 110.480 92.850 111.320 92.970 ;
        RECT 110.480 92.620 111.340 92.850 ;
        RECT 110.485 91.090 110.675 92.620 ;
        RECT 111.110 91.095 111.340 92.620 ;
        RECT 111.700 91.105 111.930 92.850 ;
        RECT 111.110 91.090 111.435 91.095 ;
        RECT 110.485 90.690 111.435 91.090 ;
        RECT 108.220 89.920 109.180 90.690 ;
        RECT 97.220 89.510 98.170 89.515 ;
        RECT 95.790 87.770 96.390 88.370 ;
        RECT 97.220 87.990 97.415 89.510 ;
        RECT 97.850 87.990 98.080 89.510 ;
        RECT 104.180 89.135 104.510 89.540 ;
        RECT 104.780 89.135 105.110 89.540 ;
        RECT 105.380 89.135 105.710 89.540 ;
        RECT 105.980 89.135 106.310 89.540 ;
        RECT 107.855 89.520 108.170 89.760 ;
        RECT 95.970 87.760 96.200 87.770 ;
        RECT 97.220 87.600 98.080 87.990 ;
        RECT 102.855 88.885 106.310 89.135 ;
        RECT 93.060 87.370 98.080 87.600 ;
        RECT 89.320 86.820 92.535 87.050 ;
        RECT 89.320 86.815 90.280 86.820 ;
        RECT 91.200 86.815 92.535 86.820 ;
        RECT 93.080 86.815 94.040 87.045 ;
        RECT 94.960 87.010 95.920 87.045 ;
        RECT 94.960 86.815 96.170 87.010 ;
        RECT 88.940 86.600 89.270 86.610 ;
        RECT 88.450 82.845 88.680 86.365 ;
        RECT 88.940 86.000 89.550 86.600 ;
        RECT 89.040 82.845 89.270 86.000 ;
        RECT 88.450 82.610 88.765 82.845 ;
        RECT 87.440 82.175 88.400 82.405 ;
        RECT 86.715 81.930 87.265 82.120 ;
        RECT 85.560 81.635 86.520 81.865 ;
        RECT 85.195 81.190 85.510 81.430 ;
        RECT 71.430 77.430 71.660 81.190 ;
        RECT 72.685 77.660 72.875 81.190 ;
        RECT 73.310 81.185 73.625 81.190 ;
        RECT 73.310 77.660 73.540 81.185 ;
        RECT 72.680 77.225 73.540 77.660 ;
        RECT 68.540 77.000 69.630 77.210 ;
        RECT 68.540 76.900 69.500 77.000 ;
        RECT 70.420 76.995 71.380 77.225 ;
        RECT 72.300 77.000 73.540 77.225 ;
        RECT 72.300 76.995 73.260 77.000 ;
        RECT 74.040 76.430 75.230 78.590 ;
        RECT 75.700 76.430 76.890 78.590 ;
        RECT 78.880 77.620 79.230 79.840 ;
        RECT 85.280 77.430 85.510 81.190 ;
        RECT 85.945 77.225 86.135 81.635 ;
        RECT 86.725 81.430 87.265 81.930 ;
        RECT 87.450 81.865 88.390 82.175 ;
        RECT 87.440 81.635 88.400 81.865 ;
        RECT 86.570 81.195 87.390 81.430 ;
        RECT 86.570 81.190 86.915 81.195 ;
        RECT 86.570 77.670 86.800 81.190 ;
        RECT 87.160 77.670 87.390 81.195 ;
        RECT 86.570 77.480 87.390 77.670 ;
        RECT 86.570 77.430 86.800 77.480 ;
        RECT 87.160 77.430 87.390 77.480 ;
        RECT 87.825 77.225 88.015 81.635 ;
        RECT 88.575 81.430 88.765 82.610 ;
        RECT 88.450 81.185 88.765 81.430 ;
        RECT 88.935 82.610 89.270 82.845 ;
        RECT 88.935 81.430 89.125 82.610 ;
        RECT 89.705 82.410 89.895 86.815 ;
        RECT 91.580 86.380 92.535 86.815 ;
        RECT 91.585 82.850 91.775 86.380 ;
        RECT 92.210 86.370 92.535 86.380 ;
        RECT 92.210 82.850 92.440 86.370 ;
        RECT 91.585 82.845 92.520 82.850 ;
        RECT 91.585 82.840 92.525 82.845 ;
        RECT 91.580 82.410 92.525 82.840 ;
        RECT 93.465 82.410 93.655 86.815 ;
        RECT 95.340 86.670 96.170 86.815 ;
        RECT 93.900 86.070 94.510 86.670 ;
        RECT 95.340 86.380 96.390 86.670 ;
        RECT 94.090 82.815 94.320 86.070 ;
        RECT 95.345 82.850 95.535 86.380 ;
        RECT 95.780 86.070 96.390 86.380 ;
        RECT 95.970 82.855 96.200 86.070 ;
        RECT 96.760 84.705 97.010 87.370 ;
        RECT 97.530 84.680 98.720 86.840 ;
        RECT 101.540 85.410 101.890 87.630 ;
        RECT 102.855 86.600 103.105 88.885 ;
        RECT 104.180 88.480 104.510 88.885 ;
        RECT 104.780 88.480 105.110 88.885 ;
        RECT 105.380 88.480 105.710 88.885 ;
        RECT 105.980 88.480 106.310 88.885 ;
        RECT 107.940 88.370 108.170 89.520 ;
        RECT 104.250 87.620 104.710 87.850 ;
        RECT 105.650 87.620 106.110 87.850 ;
        RECT 107.800 87.760 108.400 88.370 ;
        RECT 103.970 87.115 104.200 87.460 ;
        RECT 103.805 86.960 104.200 87.115 ;
        RECT 103.805 86.925 104.185 86.960 ;
        RECT 103.805 86.600 103.995 86.925 ;
        RECT 104.385 86.800 104.575 87.620 ;
        RECT 105.370 87.115 105.600 87.460 ;
        RECT 105.205 86.960 105.600 87.115 ;
        RECT 105.205 86.925 105.585 86.960 ;
        RECT 102.820 85.825 103.995 86.600 ;
        RECT 104.250 86.730 104.710 86.800 ;
        RECT 104.250 86.570 104.735 86.730 ;
        RECT 104.385 86.505 104.735 86.570 ;
        RECT 105.205 86.505 105.395 86.925 ;
        RECT 105.785 86.800 105.975 87.620 ;
        RECT 105.650 86.670 106.110 86.800 ;
        RECT 105.650 86.570 106.130 86.670 ;
        RECT 107.800 86.610 107.995 87.760 ;
        RECT 108.605 87.600 108.795 89.920 ;
        RECT 110.100 89.910 111.435 90.690 ;
        RECT 110.485 89.520 111.435 89.910 ;
        RECT 111.615 90.850 111.930 91.105 ;
        RECT 111.615 89.760 111.805 90.850 ;
        RECT 112.365 90.690 112.555 93.010 ;
        RECT 112.990 92.800 113.220 92.850 ;
        RECT 113.580 92.800 113.810 92.850 ;
        RECT 112.990 92.610 113.810 92.800 ;
        RECT 112.990 91.090 113.220 92.610 ;
        RECT 113.580 91.090 113.810 92.610 ;
        RECT 112.990 90.850 113.810 91.090 ;
        RECT 111.980 89.920 112.940 90.690 ;
        RECT 111.615 89.520 111.930 89.760 ;
        RECT 110.485 88.010 110.675 89.520 ;
        RECT 111.110 88.010 111.340 89.520 ;
        RECT 111.700 88.370 111.930 89.520 ;
        RECT 110.480 88.005 111.420 88.010 ;
        RECT 110.480 87.600 111.425 88.005 ;
        RECT 108.220 87.580 109.180 87.600 ;
        RECT 110.100 87.580 111.425 87.600 ;
        RECT 108.220 87.390 111.425 87.580 ;
        RECT 108.220 87.370 109.180 87.390 ;
        RECT 110.100 87.370 111.425 87.390 ;
        RECT 108.220 86.815 109.180 87.045 ;
        RECT 110.100 86.815 111.060 87.045 ;
        RECT 104.385 86.315 105.395 86.505 ;
        RECT 104.385 86.235 104.735 86.315 ;
        RECT 104.250 86.155 104.735 86.235 ;
        RECT 104.250 86.005 104.710 86.155 ;
        RECT 102.820 85.800 104.180 85.825 ;
        RECT 102.820 85.600 104.200 85.800 ;
        RECT 103.970 84.800 104.200 85.600 ;
        RECT 104.385 84.595 104.575 86.005 ;
        RECT 105.205 85.825 105.395 86.315 ;
        RECT 105.785 86.515 106.130 86.570 ;
        RECT 106.570 86.515 107.570 86.600 ;
        RECT 105.785 86.325 107.570 86.515 ;
        RECT 105.785 86.235 106.130 86.325 ;
        RECT 105.650 86.200 106.130 86.235 ;
        RECT 105.650 86.005 106.110 86.200 ;
        RECT 105.205 85.800 105.585 85.825 ;
        RECT 105.205 85.635 105.600 85.800 ;
        RECT 105.370 84.800 105.600 85.635 ;
        RECT 105.785 84.595 105.975 86.005 ;
        RECT 106.570 85.600 107.570 86.325 ;
        RECT 107.800 86.010 108.400 86.610 ;
        RECT 104.250 84.365 104.710 84.595 ;
        RECT 105.650 84.365 106.110 84.595 ;
        RECT 95.970 82.850 96.285 82.855 ;
        RECT 94.090 82.610 94.405 82.815 ;
        RECT 89.320 81.630 90.280 82.410 ;
        RECT 91.200 81.630 92.525 82.410 ;
        RECT 93.060 81.630 94.060 82.410 ;
        RECT 88.935 81.190 89.270 81.430 ;
        RECT 88.450 77.430 88.680 81.185 ;
        RECT 89.040 77.430 89.270 81.190 ;
        RECT 89.705 77.230 89.895 81.630 ;
        RECT 91.585 81.185 92.525 81.630 ;
        RECT 91.585 81.180 92.520 81.185 ;
        RECT 91.585 77.660 91.775 81.180 ;
        RECT 92.210 77.660 92.440 81.180 ;
        RECT 91.585 77.430 92.440 77.660 ;
        RECT 91.585 77.230 92.410 77.430 ;
        RECT 85.560 76.995 86.520 77.225 ;
        RECT 87.440 76.995 88.400 77.225 ;
        RECT 89.320 76.900 90.280 77.230 ;
        RECT 91.200 77.210 92.410 77.230 ;
        RECT 93.465 77.225 93.655 81.630 ;
        RECT 94.215 81.430 94.405 82.610 ;
        RECT 95.345 82.410 96.285 82.850 ;
        RECT 94.940 81.630 96.285 82.410 ;
        RECT 101.540 82.120 101.890 84.340 ;
        RECT 107.940 82.855 108.170 86.010 ;
        RECT 107.855 82.610 108.170 82.855 ;
        RECT 94.090 81.190 94.405 81.430 ;
        RECT 95.345 81.190 96.285 81.630 ;
        RECT 107.855 81.430 108.045 82.610 ;
        RECT 108.605 82.405 108.795 86.815 ;
        RECT 109.230 86.560 109.460 86.610 ;
        RECT 109.820 86.560 110.050 86.610 ;
        RECT 109.230 86.370 110.050 86.560 ;
        RECT 109.230 82.855 109.460 86.370 ;
        RECT 109.230 82.850 109.575 82.855 ;
        RECT 109.820 82.850 110.050 86.370 ;
        RECT 109.230 82.610 110.050 82.850 ;
        RECT 108.220 82.175 109.180 82.405 ;
        RECT 108.280 81.865 109.120 82.175 ;
        RECT 109.385 82.120 109.925 82.610 ;
        RECT 110.485 82.405 110.675 86.815 ;
        RECT 111.235 86.610 111.425 87.370 ;
        RECT 111.110 86.365 111.425 86.610 ;
        RECT 111.600 87.770 112.210 88.370 ;
        RECT 111.600 87.760 111.930 87.770 ;
        RECT 111.600 86.610 111.790 87.760 ;
        RECT 112.365 87.600 112.555 89.920 ;
        RECT 113.125 89.760 113.685 90.850 ;
        RECT 114.245 90.690 114.435 93.010 ;
        RECT 114.870 91.090 115.100 92.850 ;
        RECT 114.870 90.850 115.185 91.090 ;
        RECT 113.860 89.920 114.820 90.690 ;
        RECT 112.990 89.520 113.810 89.760 ;
        RECT 112.990 88.000 113.220 89.520 ;
        RECT 113.580 88.000 113.810 89.520 ;
        RECT 112.990 87.810 113.810 88.000 ;
        RECT 112.990 87.760 113.220 87.810 ;
        RECT 113.580 87.760 113.810 87.810 ;
        RECT 114.245 87.600 114.435 89.920 ;
        RECT 114.995 89.760 115.185 90.850 ;
        RECT 116.125 90.690 116.315 93.010 ;
        RECT 116.750 91.095 116.980 92.850 ;
        RECT 116.750 90.850 117.065 91.095 ;
        RECT 115.720 89.920 116.720 90.690 ;
        RECT 114.870 89.515 115.185 89.760 ;
        RECT 114.870 88.005 115.100 89.515 ;
        RECT 114.870 87.760 115.195 88.005 ;
        RECT 111.980 87.370 112.940 87.600 ;
        RECT 113.860 87.370 114.820 87.600 ;
        RECT 115.005 87.050 115.195 87.760 ;
        RECT 116.125 87.600 116.315 89.920 ;
        RECT 116.875 89.760 117.065 90.850 ;
        RECT 118.005 90.690 118.195 93.010 ;
        RECT 118.630 91.105 118.860 92.850 ;
        RECT 119.880 92.610 120.740 93.010 ;
        RECT 118.630 90.850 118.945 91.105 ;
        RECT 117.600 89.920 118.600 90.690 ;
        RECT 116.750 89.515 117.065 89.760 ;
        RECT 116.750 88.370 116.980 89.515 ;
        RECT 116.570 87.770 117.170 88.370 ;
        RECT 116.750 87.760 116.980 87.770 ;
        RECT 118.005 87.600 118.195 89.920 ;
        RECT 118.755 89.760 118.945 90.850 ;
        RECT 119.880 91.080 120.075 92.610 ;
        RECT 120.510 91.090 120.740 92.610 ;
        RECT 120.510 91.080 120.835 91.090 ;
        RECT 119.880 90.690 120.835 91.080 ;
        RECT 119.480 89.920 120.835 90.690 ;
        RECT 121.390 90.355 122.040 90.540 ;
        RECT 122.990 90.355 123.310 90.390 ;
        RECT 121.390 90.165 123.310 90.355 ;
        RECT 121.390 89.990 122.040 90.165 ;
        RECT 122.990 90.130 123.310 90.165 ;
        RECT 118.630 89.520 118.945 89.760 ;
        RECT 118.630 88.370 118.860 89.520 ;
        RECT 119.880 89.515 120.835 89.920 ;
        RECT 124.200 89.910 124.550 92.130 ;
        RECT 119.880 89.510 120.830 89.515 ;
        RECT 118.450 87.770 119.050 88.370 ;
        RECT 119.880 87.990 120.075 89.510 ;
        RECT 120.510 87.990 120.740 89.510 ;
        RECT 118.630 87.760 118.860 87.770 ;
        RECT 119.880 87.600 120.740 87.990 ;
        RECT 115.720 87.370 120.740 87.600 ;
        RECT 111.980 86.820 115.195 87.050 ;
        RECT 111.980 86.815 112.940 86.820 ;
        RECT 113.860 86.815 115.195 86.820 ;
        RECT 115.740 86.815 116.700 87.045 ;
        RECT 117.620 87.010 118.580 87.045 ;
        RECT 117.620 86.815 118.830 87.010 ;
        RECT 111.600 86.600 111.930 86.610 ;
        RECT 111.110 82.845 111.340 86.365 ;
        RECT 111.600 86.000 112.210 86.600 ;
        RECT 111.700 82.845 111.930 86.000 ;
        RECT 111.110 82.610 111.425 82.845 ;
        RECT 110.100 82.175 111.060 82.405 ;
        RECT 109.375 81.930 109.925 82.120 ;
        RECT 108.220 81.635 109.180 81.865 ;
        RECT 107.855 81.190 108.170 81.430 ;
        RECT 94.090 77.430 94.320 81.190 ;
        RECT 95.345 77.660 95.535 81.190 ;
        RECT 95.970 81.185 96.285 81.190 ;
        RECT 95.970 77.660 96.200 81.185 ;
        RECT 95.340 77.225 96.200 77.660 ;
        RECT 91.200 77.000 92.290 77.210 ;
        RECT 91.200 76.900 92.160 77.000 ;
        RECT 93.080 76.995 94.040 77.225 ;
        RECT 94.960 77.000 96.200 77.225 ;
        RECT 94.960 76.995 95.920 77.000 ;
        RECT 96.700 76.430 97.890 78.590 ;
        RECT 98.360 76.430 99.550 78.590 ;
        RECT 101.540 77.620 101.890 79.840 ;
        RECT 107.940 77.430 108.170 81.190 ;
        RECT 108.605 77.225 108.795 81.635 ;
        RECT 109.385 81.430 109.925 81.930 ;
        RECT 110.110 81.865 111.050 82.175 ;
        RECT 110.100 81.635 111.060 81.865 ;
        RECT 109.230 81.195 110.050 81.430 ;
        RECT 109.230 81.190 109.575 81.195 ;
        RECT 109.230 77.670 109.460 81.190 ;
        RECT 109.820 77.670 110.050 81.195 ;
        RECT 109.230 77.480 110.050 77.670 ;
        RECT 109.230 77.430 109.460 77.480 ;
        RECT 109.820 77.430 110.050 77.480 ;
        RECT 110.485 77.225 110.675 81.635 ;
        RECT 111.235 81.430 111.425 82.610 ;
        RECT 111.110 81.185 111.425 81.430 ;
        RECT 111.595 82.610 111.930 82.845 ;
        RECT 111.595 81.430 111.785 82.610 ;
        RECT 112.365 82.410 112.555 86.815 ;
        RECT 114.240 86.380 115.195 86.815 ;
        RECT 114.245 82.850 114.435 86.380 ;
        RECT 114.870 86.370 115.195 86.380 ;
        RECT 114.870 82.850 115.100 86.370 ;
        RECT 114.245 82.845 115.180 82.850 ;
        RECT 114.245 82.840 115.185 82.845 ;
        RECT 114.240 82.410 115.185 82.840 ;
        RECT 116.125 82.410 116.315 86.815 ;
        RECT 118.000 86.670 118.830 86.815 ;
        RECT 116.560 86.070 117.170 86.670 ;
        RECT 118.000 86.380 119.050 86.670 ;
        RECT 116.750 82.815 116.980 86.070 ;
        RECT 118.005 82.850 118.195 86.380 ;
        RECT 118.440 86.070 119.050 86.380 ;
        RECT 118.630 82.855 118.860 86.070 ;
        RECT 119.420 84.705 119.670 87.370 ;
        RECT 120.190 84.680 121.380 86.840 ;
        RECT 124.200 85.410 124.550 87.630 ;
        RECT 118.630 82.850 118.945 82.855 ;
        RECT 116.750 82.610 117.065 82.815 ;
        RECT 111.980 81.630 112.940 82.410 ;
        RECT 113.860 81.630 115.185 82.410 ;
        RECT 115.720 81.630 116.720 82.410 ;
        RECT 111.595 81.190 111.930 81.430 ;
        RECT 111.110 77.430 111.340 81.185 ;
        RECT 111.700 77.430 111.930 81.190 ;
        RECT 112.365 77.230 112.555 81.630 ;
        RECT 114.245 81.185 115.185 81.630 ;
        RECT 114.245 81.180 115.180 81.185 ;
        RECT 114.245 77.660 114.435 81.180 ;
        RECT 114.870 77.660 115.100 81.180 ;
        RECT 114.245 77.430 115.100 77.660 ;
        RECT 114.245 77.230 115.070 77.430 ;
        RECT 108.220 76.995 109.180 77.225 ;
        RECT 110.100 76.995 111.060 77.225 ;
        RECT 111.980 76.900 112.940 77.230 ;
        RECT 113.860 77.210 115.070 77.230 ;
        RECT 116.125 77.225 116.315 81.630 ;
        RECT 116.875 81.430 117.065 82.610 ;
        RECT 118.005 82.410 118.945 82.850 ;
        RECT 117.600 81.630 118.945 82.410 ;
        RECT 124.200 82.120 124.550 84.340 ;
        RECT 116.750 81.190 117.065 81.430 ;
        RECT 118.005 81.190 118.945 81.630 ;
        RECT 116.750 77.430 116.980 81.190 ;
        RECT 118.005 77.660 118.195 81.190 ;
        RECT 118.630 81.185 118.945 81.190 ;
        RECT 118.630 77.660 118.860 81.185 ;
        RECT 118.000 77.225 118.860 77.660 ;
        RECT 113.860 77.000 114.950 77.210 ;
        RECT 113.860 76.900 114.820 77.000 ;
        RECT 115.740 76.995 116.700 77.225 ;
        RECT 117.620 77.000 118.860 77.225 ;
        RECT 117.620 76.995 118.580 77.000 ;
        RECT 119.360 76.430 120.550 78.590 ;
        RECT 121.020 76.430 122.210 78.590 ;
        RECT 124.200 77.620 124.550 79.840 ;
        RECT 40.270 75.900 41.170 75.950 ;
        RECT 42.150 75.900 43.050 75.950 ;
        RECT 40.240 75.670 41.200 75.900 ;
        RECT 42.120 75.875 43.080 75.900 ;
        RECT 42.120 75.670 43.340 75.875 ;
        RECT 44.000 75.670 44.960 75.900 ;
        RECT 45.880 75.670 46.840 75.900 ;
        RECT 47.740 75.670 48.740 75.990 ;
        RECT 49.620 75.670 50.620 75.990 ;
        RECT 51.500 75.900 52.500 75.990 ;
        RECT 62.930 75.900 63.830 75.950 ;
        RECT 64.810 75.900 65.710 75.950 ;
        RECT 51.500 75.670 52.760 75.900 ;
        RECT 62.900 75.670 63.860 75.900 ;
        RECT 64.780 75.875 65.740 75.900 ;
        RECT 64.780 75.670 66.000 75.875 ;
        RECT 66.660 75.670 67.620 75.900 ;
        RECT 68.540 75.670 69.500 75.900 ;
        RECT 70.400 75.670 71.400 75.990 ;
        RECT 72.280 75.670 73.280 75.990 ;
        RECT 74.160 75.900 75.160 75.990 ;
        RECT 85.590 75.900 86.490 75.950 ;
        RECT 87.470 75.900 88.370 75.950 ;
        RECT 74.160 75.670 75.420 75.900 ;
        RECT 85.560 75.670 86.520 75.900 ;
        RECT 87.440 75.875 88.400 75.900 ;
        RECT 87.440 75.670 88.660 75.875 ;
        RECT 89.320 75.670 90.280 75.900 ;
        RECT 91.200 75.670 92.160 75.900 ;
        RECT 93.060 75.670 94.060 75.990 ;
        RECT 94.940 75.670 95.940 75.990 ;
        RECT 96.820 75.900 97.820 75.990 ;
        RECT 108.250 75.900 109.150 75.950 ;
        RECT 110.130 75.900 111.030 75.950 ;
        RECT 96.820 75.670 98.080 75.900 ;
        RECT 108.220 75.670 109.180 75.900 ;
        RECT 110.100 75.875 111.060 75.900 ;
        RECT 110.100 75.670 111.320 75.875 ;
        RECT 111.980 75.670 112.940 75.900 ;
        RECT 113.860 75.670 114.820 75.900 ;
        RECT 115.720 75.670 116.720 75.990 ;
        RECT 117.600 75.670 118.600 75.990 ;
        RECT 119.480 75.900 120.480 75.990 ;
        RECT 119.480 75.670 120.740 75.900 ;
        RECT 40.270 75.630 41.170 75.670 ;
        RECT 42.150 75.630 43.340 75.670 ;
        RECT 39.960 73.745 40.190 75.510 ;
        RECT 39.875 73.510 40.190 73.745 ;
        RECT 39.875 72.420 40.065 73.510 ;
        RECT 40.625 73.350 40.815 75.630 ;
        RECT 42.500 75.510 43.340 75.630 ;
        RECT 42.500 75.280 43.360 75.510 ;
        RECT 42.505 73.750 42.695 75.280 ;
        RECT 43.130 73.755 43.360 75.280 ;
        RECT 43.720 73.765 43.950 75.510 ;
        RECT 43.130 73.750 43.455 73.755 ;
        RECT 42.505 73.350 43.455 73.750 ;
        RECT 40.240 72.580 41.200 73.350 ;
        RECT 36.200 71.795 36.530 72.200 ;
        RECT 36.800 71.795 37.130 72.200 ;
        RECT 37.400 71.795 37.730 72.200 ;
        RECT 38.000 71.795 38.330 72.200 ;
        RECT 39.875 72.180 40.190 72.420 ;
        RECT 34.875 71.545 38.330 71.795 ;
        RECT 34.875 69.260 35.125 71.545 ;
        RECT 36.200 71.140 36.530 71.545 ;
        RECT 36.800 71.140 37.130 71.545 ;
        RECT 37.400 71.140 37.730 71.545 ;
        RECT 38.000 71.140 38.330 71.545 ;
        RECT 39.960 71.030 40.190 72.180 ;
        RECT 36.270 70.280 36.730 70.510 ;
        RECT 37.670 70.280 38.130 70.510 ;
        RECT 39.820 70.420 40.420 71.030 ;
        RECT 35.990 69.775 36.220 70.120 ;
        RECT 35.825 69.620 36.220 69.775 ;
        RECT 35.825 69.585 36.205 69.620 ;
        RECT 35.825 69.260 36.015 69.585 ;
        RECT 36.405 69.460 36.595 70.280 ;
        RECT 37.390 69.775 37.620 70.120 ;
        RECT 37.225 69.620 37.620 69.775 ;
        RECT 37.225 69.585 37.605 69.620 ;
        RECT 34.840 68.485 36.015 69.260 ;
        RECT 36.270 69.390 36.730 69.460 ;
        RECT 36.270 69.230 36.755 69.390 ;
        RECT 36.405 69.165 36.755 69.230 ;
        RECT 37.225 69.165 37.415 69.585 ;
        RECT 37.805 69.460 37.995 70.280 ;
        RECT 37.670 69.330 38.130 69.460 ;
        RECT 37.670 69.230 38.150 69.330 ;
        RECT 39.820 69.270 40.015 70.420 ;
        RECT 40.625 70.260 40.815 72.580 ;
        RECT 42.120 72.570 43.455 73.350 ;
        RECT 42.505 72.180 43.455 72.570 ;
        RECT 43.635 73.510 43.950 73.765 ;
        RECT 43.635 72.420 43.825 73.510 ;
        RECT 44.385 73.350 44.575 75.670 ;
        RECT 45.010 75.460 45.240 75.510 ;
        RECT 45.600 75.460 45.830 75.510 ;
        RECT 45.010 75.270 45.830 75.460 ;
        RECT 45.010 73.750 45.240 75.270 ;
        RECT 45.600 73.750 45.830 75.270 ;
        RECT 45.010 73.510 45.830 73.750 ;
        RECT 44.000 72.580 44.960 73.350 ;
        RECT 43.635 72.180 43.950 72.420 ;
        RECT 42.505 70.670 42.695 72.180 ;
        RECT 43.130 70.670 43.360 72.180 ;
        RECT 43.720 71.030 43.950 72.180 ;
        RECT 42.500 70.665 43.440 70.670 ;
        RECT 42.500 70.260 43.445 70.665 ;
        RECT 40.240 70.240 41.200 70.260 ;
        RECT 42.120 70.240 43.445 70.260 ;
        RECT 40.240 70.050 43.445 70.240 ;
        RECT 40.240 70.030 41.200 70.050 ;
        RECT 42.120 70.030 43.445 70.050 ;
        RECT 40.240 69.475 41.200 69.705 ;
        RECT 42.120 69.475 43.080 69.705 ;
        RECT 36.405 68.975 37.415 69.165 ;
        RECT 36.405 68.895 36.755 68.975 ;
        RECT 36.270 68.815 36.755 68.895 ;
        RECT 36.270 68.665 36.730 68.815 ;
        RECT 34.840 68.460 36.200 68.485 ;
        RECT 34.840 68.260 36.220 68.460 ;
        RECT 35.990 67.460 36.220 68.260 ;
        RECT 36.405 67.255 36.595 68.665 ;
        RECT 37.225 68.485 37.415 68.975 ;
        RECT 37.805 69.175 38.150 69.230 ;
        RECT 38.590 69.175 39.590 69.260 ;
        RECT 37.805 68.985 39.590 69.175 ;
        RECT 37.805 68.895 38.150 68.985 ;
        RECT 37.670 68.860 38.150 68.895 ;
        RECT 37.670 68.665 38.130 68.860 ;
        RECT 37.225 68.460 37.605 68.485 ;
        RECT 37.225 68.295 37.620 68.460 ;
        RECT 37.390 67.460 37.620 68.295 ;
        RECT 37.805 67.255 37.995 68.665 ;
        RECT 38.590 68.260 39.590 68.985 ;
        RECT 39.820 68.670 40.420 69.270 ;
        RECT 36.270 67.025 36.730 67.255 ;
        RECT 37.670 67.025 38.130 67.255 ;
        RECT 39.960 65.515 40.190 68.670 ;
        RECT 39.875 65.270 40.190 65.515 ;
        RECT 39.875 64.090 40.065 65.270 ;
        RECT 40.625 65.065 40.815 69.475 ;
        RECT 41.250 69.220 41.480 69.270 ;
        RECT 41.840 69.220 42.070 69.270 ;
        RECT 41.250 69.030 42.070 69.220 ;
        RECT 41.250 65.515 41.480 69.030 ;
        RECT 41.250 65.510 41.595 65.515 ;
        RECT 41.840 65.510 42.070 69.030 ;
        RECT 41.250 65.270 42.070 65.510 ;
        RECT 40.240 64.835 41.200 65.065 ;
        RECT 40.300 64.525 41.140 64.835 ;
        RECT 41.405 64.780 41.945 65.270 ;
        RECT 42.505 65.065 42.695 69.475 ;
        RECT 43.255 69.270 43.445 70.030 ;
        RECT 43.130 69.025 43.445 69.270 ;
        RECT 43.620 70.430 44.230 71.030 ;
        RECT 43.620 70.420 43.950 70.430 ;
        RECT 43.620 69.270 43.810 70.420 ;
        RECT 44.385 70.260 44.575 72.580 ;
        RECT 45.145 72.420 45.705 73.510 ;
        RECT 46.265 73.350 46.455 75.670 ;
        RECT 46.890 73.750 47.120 75.510 ;
        RECT 46.890 73.510 47.205 73.750 ;
        RECT 45.880 72.580 46.840 73.350 ;
        RECT 45.010 72.180 45.830 72.420 ;
        RECT 45.010 70.660 45.240 72.180 ;
        RECT 45.600 70.660 45.830 72.180 ;
        RECT 45.010 70.470 45.830 70.660 ;
        RECT 45.010 70.420 45.240 70.470 ;
        RECT 45.600 70.420 45.830 70.470 ;
        RECT 46.265 70.260 46.455 72.580 ;
        RECT 47.015 72.420 47.205 73.510 ;
        RECT 48.145 73.350 48.335 75.670 ;
        RECT 48.770 73.755 49.000 75.510 ;
        RECT 48.770 73.510 49.085 73.755 ;
        RECT 47.740 72.580 48.740 73.350 ;
        RECT 46.890 72.175 47.205 72.420 ;
        RECT 46.890 70.665 47.120 72.175 ;
        RECT 46.890 70.420 47.215 70.665 ;
        RECT 44.000 70.030 44.960 70.260 ;
        RECT 45.880 70.030 46.840 70.260 ;
        RECT 47.025 69.710 47.215 70.420 ;
        RECT 48.145 70.260 48.335 72.580 ;
        RECT 48.895 72.420 49.085 73.510 ;
        RECT 50.025 73.350 50.215 75.670 ;
        RECT 50.650 73.765 50.880 75.510 ;
        RECT 51.900 75.270 52.760 75.670 ;
        RECT 62.930 75.630 63.830 75.670 ;
        RECT 64.810 75.630 66.000 75.670 ;
        RECT 50.650 73.510 50.965 73.765 ;
        RECT 49.620 72.580 50.620 73.350 ;
        RECT 48.770 72.175 49.085 72.420 ;
        RECT 48.770 71.030 49.000 72.175 ;
        RECT 48.590 70.430 49.190 71.030 ;
        RECT 48.770 70.420 49.000 70.430 ;
        RECT 50.025 70.260 50.215 72.580 ;
        RECT 50.775 72.420 50.965 73.510 ;
        RECT 51.900 73.740 52.095 75.270 ;
        RECT 52.530 73.750 52.760 75.270 ;
        RECT 52.530 73.740 52.855 73.750 ;
        RECT 51.900 73.350 52.855 73.740 ;
        RECT 51.500 72.580 52.855 73.350 ;
        RECT 53.410 73.015 54.060 73.200 ;
        RECT 55.010 73.015 55.330 73.050 ;
        RECT 53.410 72.825 55.330 73.015 ;
        RECT 53.410 72.650 54.060 72.825 ;
        RECT 55.010 72.790 55.330 72.825 ;
        RECT 50.650 72.180 50.965 72.420 ;
        RECT 50.650 71.030 50.880 72.180 ;
        RECT 51.900 72.175 52.855 72.580 ;
        RECT 56.220 72.570 56.570 74.790 ;
        RECT 62.620 73.745 62.850 75.510 ;
        RECT 62.535 73.510 62.850 73.745 ;
        RECT 62.535 72.420 62.725 73.510 ;
        RECT 63.285 73.350 63.475 75.630 ;
        RECT 65.160 75.510 66.000 75.630 ;
        RECT 65.160 75.280 66.020 75.510 ;
        RECT 65.165 73.750 65.355 75.280 ;
        RECT 65.790 73.755 66.020 75.280 ;
        RECT 66.380 73.765 66.610 75.510 ;
        RECT 65.790 73.750 66.115 73.755 ;
        RECT 65.165 73.350 66.115 73.750 ;
        RECT 62.900 72.580 63.860 73.350 ;
        RECT 51.900 72.170 52.850 72.175 ;
        RECT 50.470 70.430 51.070 71.030 ;
        RECT 51.900 70.650 52.095 72.170 ;
        RECT 52.530 70.650 52.760 72.170 ;
        RECT 58.860 71.795 59.190 72.200 ;
        RECT 59.460 71.795 59.790 72.200 ;
        RECT 60.060 71.795 60.390 72.200 ;
        RECT 60.660 71.795 60.990 72.200 ;
        RECT 62.535 72.180 62.850 72.420 ;
        RECT 50.650 70.420 50.880 70.430 ;
        RECT 51.900 70.260 52.760 70.650 ;
        RECT 57.535 71.545 60.990 71.795 ;
        RECT 47.740 70.030 52.760 70.260 ;
        RECT 44.000 69.480 47.215 69.710 ;
        RECT 44.000 69.475 44.960 69.480 ;
        RECT 45.880 69.475 47.215 69.480 ;
        RECT 47.760 69.475 48.720 69.705 ;
        RECT 49.640 69.670 50.600 69.705 ;
        RECT 49.640 69.475 50.850 69.670 ;
        RECT 43.620 69.260 43.950 69.270 ;
        RECT 43.130 65.505 43.360 69.025 ;
        RECT 43.620 68.660 44.230 69.260 ;
        RECT 43.720 65.505 43.950 68.660 ;
        RECT 43.130 65.270 43.445 65.505 ;
        RECT 42.120 64.835 43.080 65.065 ;
        RECT 41.395 64.590 41.945 64.780 ;
        RECT 40.240 64.295 41.200 64.525 ;
        RECT 39.875 63.850 40.190 64.090 ;
        RECT 39.960 60.090 40.190 63.850 ;
        RECT 40.625 59.885 40.815 64.295 ;
        RECT 41.405 64.090 41.945 64.590 ;
        RECT 42.130 64.525 43.070 64.835 ;
        RECT 42.120 64.295 43.080 64.525 ;
        RECT 41.250 63.855 42.070 64.090 ;
        RECT 41.250 63.850 41.595 63.855 ;
        RECT 41.250 60.330 41.480 63.850 ;
        RECT 41.840 60.330 42.070 63.855 ;
        RECT 41.250 60.140 42.070 60.330 ;
        RECT 41.250 60.090 41.480 60.140 ;
        RECT 41.840 60.090 42.070 60.140 ;
        RECT 42.505 59.885 42.695 64.295 ;
        RECT 43.255 64.090 43.445 65.270 ;
        RECT 43.130 63.845 43.445 64.090 ;
        RECT 43.615 65.270 43.950 65.505 ;
        RECT 43.615 64.090 43.805 65.270 ;
        RECT 44.385 65.070 44.575 69.475 ;
        RECT 46.260 69.040 47.215 69.475 ;
        RECT 46.265 65.510 46.455 69.040 ;
        RECT 46.890 69.030 47.215 69.040 ;
        RECT 46.890 65.510 47.120 69.030 ;
        RECT 46.265 65.505 47.200 65.510 ;
        RECT 46.265 65.500 47.205 65.505 ;
        RECT 46.260 65.070 47.205 65.500 ;
        RECT 48.145 65.070 48.335 69.475 ;
        RECT 50.020 69.330 50.850 69.475 ;
        RECT 48.580 68.730 49.190 69.330 ;
        RECT 50.020 69.040 51.070 69.330 ;
        RECT 48.770 65.475 49.000 68.730 ;
        RECT 50.025 65.510 50.215 69.040 ;
        RECT 50.460 68.730 51.070 69.040 ;
        RECT 50.650 65.515 50.880 68.730 ;
        RECT 51.440 67.365 51.690 70.030 ;
        RECT 52.210 67.340 53.400 69.500 ;
        RECT 56.220 68.070 56.570 70.290 ;
        RECT 57.535 69.260 57.785 71.545 ;
        RECT 58.860 71.140 59.190 71.545 ;
        RECT 59.460 71.140 59.790 71.545 ;
        RECT 60.060 71.140 60.390 71.545 ;
        RECT 60.660 71.140 60.990 71.545 ;
        RECT 62.620 71.030 62.850 72.180 ;
        RECT 58.930 70.280 59.390 70.510 ;
        RECT 60.330 70.280 60.790 70.510 ;
        RECT 62.480 70.420 63.080 71.030 ;
        RECT 58.650 69.775 58.880 70.120 ;
        RECT 58.485 69.620 58.880 69.775 ;
        RECT 58.485 69.585 58.865 69.620 ;
        RECT 58.485 69.260 58.675 69.585 ;
        RECT 59.065 69.460 59.255 70.280 ;
        RECT 60.050 69.775 60.280 70.120 ;
        RECT 59.885 69.620 60.280 69.775 ;
        RECT 59.885 69.585 60.265 69.620 ;
        RECT 57.500 68.485 58.675 69.260 ;
        RECT 58.930 69.390 59.390 69.460 ;
        RECT 58.930 69.230 59.415 69.390 ;
        RECT 59.065 69.165 59.415 69.230 ;
        RECT 59.885 69.165 60.075 69.585 ;
        RECT 60.465 69.460 60.655 70.280 ;
        RECT 60.330 69.330 60.790 69.460 ;
        RECT 60.330 69.230 60.810 69.330 ;
        RECT 62.480 69.270 62.675 70.420 ;
        RECT 63.285 70.260 63.475 72.580 ;
        RECT 64.780 72.570 66.115 73.350 ;
        RECT 65.165 72.180 66.115 72.570 ;
        RECT 66.295 73.510 66.610 73.765 ;
        RECT 66.295 72.420 66.485 73.510 ;
        RECT 67.045 73.350 67.235 75.670 ;
        RECT 67.670 75.460 67.900 75.510 ;
        RECT 68.260 75.460 68.490 75.510 ;
        RECT 67.670 75.270 68.490 75.460 ;
        RECT 67.670 73.750 67.900 75.270 ;
        RECT 68.260 73.750 68.490 75.270 ;
        RECT 67.670 73.510 68.490 73.750 ;
        RECT 66.660 72.580 67.620 73.350 ;
        RECT 66.295 72.180 66.610 72.420 ;
        RECT 65.165 70.670 65.355 72.180 ;
        RECT 65.790 70.670 66.020 72.180 ;
        RECT 66.380 71.030 66.610 72.180 ;
        RECT 65.160 70.665 66.100 70.670 ;
        RECT 65.160 70.260 66.105 70.665 ;
        RECT 62.900 70.240 63.860 70.260 ;
        RECT 64.780 70.240 66.105 70.260 ;
        RECT 62.900 70.050 66.105 70.240 ;
        RECT 62.900 70.030 63.860 70.050 ;
        RECT 64.780 70.030 66.105 70.050 ;
        RECT 62.900 69.475 63.860 69.705 ;
        RECT 64.780 69.475 65.740 69.705 ;
        RECT 59.065 68.975 60.075 69.165 ;
        RECT 59.065 68.895 59.415 68.975 ;
        RECT 58.930 68.815 59.415 68.895 ;
        RECT 58.930 68.665 59.390 68.815 ;
        RECT 57.500 68.460 58.860 68.485 ;
        RECT 57.500 68.260 58.880 68.460 ;
        RECT 58.650 67.460 58.880 68.260 ;
        RECT 59.065 67.255 59.255 68.665 ;
        RECT 59.885 68.485 60.075 68.975 ;
        RECT 60.465 69.175 60.810 69.230 ;
        RECT 61.250 69.175 62.250 69.260 ;
        RECT 60.465 68.985 62.250 69.175 ;
        RECT 60.465 68.895 60.810 68.985 ;
        RECT 60.330 68.860 60.810 68.895 ;
        RECT 60.330 68.665 60.790 68.860 ;
        RECT 59.885 68.460 60.265 68.485 ;
        RECT 59.885 68.295 60.280 68.460 ;
        RECT 60.050 67.460 60.280 68.295 ;
        RECT 60.465 67.255 60.655 68.665 ;
        RECT 61.250 68.260 62.250 68.985 ;
        RECT 62.480 68.670 63.080 69.270 ;
        RECT 58.930 67.025 59.390 67.255 ;
        RECT 60.330 67.025 60.790 67.255 ;
        RECT 50.650 65.510 50.965 65.515 ;
        RECT 48.770 65.270 49.085 65.475 ;
        RECT 44.000 64.290 44.960 65.070 ;
        RECT 45.880 64.290 47.205 65.070 ;
        RECT 47.740 64.290 48.740 65.070 ;
        RECT 43.615 63.850 43.950 64.090 ;
        RECT 43.130 60.090 43.360 63.845 ;
        RECT 43.720 60.090 43.950 63.850 ;
        RECT 44.385 59.890 44.575 64.290 ;
        RECT 46.265 63.845 47.205 64.290 ;
        RECT 46.265 63.840 47.200 63.845 ;
        RECT 46.265 60.320 46.455 63.840 ;
        RECT 46.890 60.320 47.120 63.840 ;
        RECT 46.265 60.090 47.120 60.320 ;
        RECT 46.265 59.890 47.090 60.090 ;
        RECT 40.240 59.655 41.200 59.885 ;
        RECT 42.120 59.655 43.080 59.885 ;
        RECT 44.000 59.560 44.960 59.890 ;
        RECT 45.880 59.870 47.090 59.890 ;
        RECT 48.145 59.885 48.335 64.290 ;
        RECT 48.895 64.090 49.085 65.270 ;
        RECT 50.025 65.070 50.965 65.510 ;
        RECT 49.620 64.290 50.965 65.070 ;
        RECT 56.220 64.780 56.570 67.000 ;
        RECT 62.620 65.515 62.850 68.670 ;
        RECT 62.535 65.270 62.850 65.515 ;
        RECT 48.770 63.850 49.085 64.090 ;
        RECT 50.025 63.850 50.965 64.290 ;
        RECT 62.535 64.090 62.725 65.270 ;
        RECT 63.285 65.065 63.475 69.475 ;
        RECT 63.910 69.220 64.140 69.270 ;
        RECT 64.500 69.220 64.730 69.270 ;
        RECT 63.910 69.030 64.730 69.220 ;
        RECT 63.910 65.515 64.140 69.030 ;
        RECT 63.910 65.510 64.255 65.515 ;
        RECT 64.500 65.510 64.730 69.030 ;
        RECT 63.910 65.270 64.730 65.510 ;
        RECT 62.900 64.835 63.860 65.065 ;
        RECT 62.960 64.525 63.800 64.835 ;
        RECT 64.065 64.780 64.605 65.270 ;
        RECT 65.165 65.065 65.355 69.475 ;
        RECT 65.915 69.270 66.105 70.030 ;
        RECT 65.790 69.025 66.105 69.270 ;
        RECT 66.280 70.430 66.890 71.030 ;
        RECT 66.280 70.420 66.610 70.430 ;
        RECT 66.280 69.270 66.470 70.420 ;
        RECT 67.045 70.260 67.235 72.580 ;
        RECT 67.805 72.420 68.365 73.510 ;
        RECT 68.925 73.350 69.115 75.670 ;
        RECT 69.550 73.750 69.780 75.510 ;
        RECT 69.550 73.510 69.865 73.750 ;
        RECT 68.540 72.580 69.500 73.350 ;
        RECT 67.670 72.180 68.490 72.420 ;
        RECT 67.670 70.660 67.900 72.180 ;
        RECT 68.260 70.660 68.490 72.180 ;
        RECT 67.670 70.470 68.490 70.660 ;
        RECT 67.670 70.420 67.900 70.470 ;
        RECT 68.260 70.420 68.490 70.470 ;
        RECT 68.925 70.260 69.115 72.580 ;
        RECT 69.675 72.420 69.865 73.510 ;
        RECT 70.805 73.350 70.995 75.670 ;
        RECT 71.430 73.755 71.660 75.510 ;
        RECT 71.430 73.510 71.745 73.755 ;
        RECT 70.400 72.580 71.400 73.350 ;
        RECT 69.550 72.175 69.865 72.420 ;
        RECT 69.550 70.665 69.780 72.175 ;
        RECT 69.550 70.420 69.875 70.665 ;
        RECT 66.660 70.030 67.620 70.260 ;
        RECT 68.540 70.030 69.500 70.260 ;
        RECT 69.685 69.710 69.875 70.420 ;
        RECT 70.805 70.260 70.995 72.580 ;
        RECT 71.555 72.420 71.745 73.510 ;
        RECT 72.685 73.350 72.875 75.670 ;
        RECT 73.310 73.765 73.540 75.510 ;
        RECT 74.560 75.270 75.420 75.670 ;
        RECT 85.590 75.630 86.490 75.670 ;
        RECT 87.470 75.630 88.660 75.670 ;
        RECT 73.310 73.510 73.625 73.765 ;
        RECT 72.280 72.580 73.280 73.350 ;
        RECT 71.430 72.175 71.745 72.420 ;
        RECT 71.430 71.030 71.660 72.175 ;
        RECT 71.250 70.430 71.850 71.030 ;
        RECT 71.430 70.420 71.660 70.430 ;
        RECT 72.685 70.260 72.875 72.580 ;
        RECT 73.435 72.420 73.625 73.510 ;
        RECT 74.560 73.740 74.755 75.270 ;
        RECT 75.190 73.750 75.420 75.270 ;
        RECT 75.190 73.740 75.515 73.750 ;
        RECT 74.560 73.350 75.515 73.740 ;
        RECT 74.160 72.580 75.515 73.350 ;
        RECT 76.070 73.015 76.720 73.200 ;
        RECT 77.670 73.015 77.990 73.050 ;
        RECT 76.070 72.825 77.990 73.015 ;
        RECT 76.070 72.650 76.720 72.825 ;
        RECT 77.670 72.790 77.990 72.825 ;
        RECT 73.310 72.180 73.625 72.420 ;
        RECT 73.310 71.030 73.540 72.180 ;
        RECT 74.560 72.175 75.515 72.580 ;
        RECT 78.880 72.570 79.230 74.790 ;
        RECT 85.280 73.745 85.510 75.510 ;
        RECT 85.195 73.510 85.510 73.745 ;
        RECT 85.195 72.420 85.385 73.510 ;
        RECT 85.945 73.350 86.135 75.630 ;
        RECT 87.820 75.510 88.660 75.630 ;
        RECT 87.820 75.280 88.680 75.510 ;
        RECT 87.825 73.750 88.015 75.280 ;
        RECT 88.450 73.755 88.680 75.280 ;
        RECT 89.040 73.765 89.270 75.510 ;
        RECT 88.450 73.750 88.775 73.755 ;
        RECT 87.825 73.350 88.775 73.750 ;
        RECT 85.560 72.580 86.520 73.350 ;
        RECT 74.560 72.170 75.510 72.175 ;
        RECT 73.130 70.430 73.730 71.030 ;
        RECT 74.560 70.650 74.755 72.170 ;
        RECT 75.190 70.650 75.420 72.170 ;
        RECT 81.520 71.795 81.850 72.200 ;
        RECT 82.120 71.795 82.450 72.200 ;
        RECT 82.720 71.795 83.050 72.200 ;
        RECT 83.320 71.795 83.650 72.200 ;
        RECT 85.195 72.180 85.510 72.420 ;
        RECT 73.310 70.420 73.540 70.430 ;
        RECT 74.560 70.260 75.420 70.650 ;
        RECT 80.195 71.545 83.650 71.795 ;
        RECT 70.400 70.030 75.420 70.260 ;
        RECT 66.660 69.480 69.875 69.710 ;
        RECT 66.660 69.475 67.620 69.480 ;
        RECT 68.540 69.475 69.875 69.480 ;
        RECT 70.420 69.475 71.380 69.705 ;
        RECT 72.300 69.670 73.260 69.705 ;
        RECT 72.300 69.475 73.510 69.670 ;
        RECT 66.280 69.260 66.610 69.270 ;
        RECT 65.790 65.505 66.020 69.025 ;
        RECT 66.280 68.660 66.890 69.260 ;
        RECT 66.380 65.505 66.610 68.660 ;
        RECT 65.790 65.270 66.105 65.505 ;
        RECT 64.780 64.835 65.740 65.065 ;
        RECT 64.055 64.590 64.605 64.780 ;
        RECT 62.900 64.295 63.860 64.525 ;
        RECT 62.535 63.850 62.850 64.090 ;
        RECT 48.770 60.090 49.000 63.850 ;
        RECT 50.025 60.320 50.215 63.850 ;
        RECT 50.650 63.845 50.965 63.850 ;
        RECT 50.650 60.320 50.880 63.845 ;
        RECT 50.020 59.885 50.880 60.320 ;
        RECT 45.880 59.660 46.970 59.870 ;
        RECT 45.880 59.560 46.840 59.660 ;
        RECT 47.760 59.655 48.720 59.885 ;
        RECT 49.640 59.660 50.880 59.885 ;
        RECT 49.640 59.655 50.600 59.660 ;
        RECT 51.380 59.090 52.570 61.250 ;
        RECT 53.040 59.090 54.230 61.250 ;
        RECT 56.220 60.280 56.570 62.500 ;
        RECT 62.620 60.090 62.850 63.850 ;
        RECT 63.285 59.885 63.475 64.295 ;
        RECT 64.065 64.090 64.605 64.590 ;
        RECT 64.790 64.525 65.730 64.835 ;
        RECT 64.780 64.295 65.740 64.525 ;
        RECT 63.910 63.855 64.730 64.090 ;
        RECT 63.910 63.850 64.255 63.855 ;
        RECT 63.910 60.330 64.140 63.850 ;
        RECT 64.500 60.330 64.730 63.855 ;
        RECT 63.910 60.140 64.730 60.330 ;
        RECT 63.910 60.090 64.140 60.140 ;
        RECT 64.500 60.090 64.730 60.140 ;
        RECT 65.165 59.885 65.355 64.295 ;
        RECT 65.915 64.090 66.105 65.270 ;
        RECT 65.790 63.845 66.105 64.090 ;
        RECT 66.275 65.270 66.610 65.505 ;
        RECT 66.275 64.090 66.465 65.270 ;
        RECT 67.045 65.070 67.235 69.475 ;
        RECT 68.920 69.040 69.875 69.475 ;
        RECT 68.925 65.510 69.115 69.040 ;
        RECT 69.550 69.030 69.875 69.040 ;
        RECT 69.550 65.510 69.780 69.030 ;
        RECT 68.925 65.505 69.860 65.510 ;
        RECT 68.925 65.500 69.865 65.505 ;
        RECT 68.920 65.070 69.865 65.500 ;
        RECT 70.805 65.070 70.995 69.475 ;
        RECT 72.680 69.330 73.510 69.475 ;
        RECT 71.240 68.730 71.850 69.330 ;
        RECT 72.680 69.040 73.730 69.330 ;
        RECT 71.430 65.475 71.660 68.730 ;
        RECT 72.685 65.510 72.875 69.040 ;
        RECT 73.120 68.730 73.730 69.040 ;
        RECT 73.310 65.515 73.540 68.730 ;
        RECT 74.100 67.365 74.350 70.030 ;
        RECT 74.870 67.340 76.060 69.500 ;
        RECT 78.880 68.070 79.230 70.290 ;
        RECT 80.195 69.260 80.445 71.545 ;
        RECT 81.520 71.140 81.850 71.545 ;
        RECT 82.120 71.140 82.450 71.545 ;
        RECT 82.720 71.140 83.050 71.545 ;
        RECT 83.320 71.140 83.650 71.545 ;
        RECT 85.280 71.030 85.510 72.180 ;
        RECT 81.590 70.280 82.050 70.510 ;
        RECT 82.990 70.280 83.450 70.510 ;
        RECT 85.140 70.420 85.740 71.030 ;
        RECT 81.310 69.775 81.540 70.120 ;
        RECT 81.145 69.620 81.540 69.775 ;
        RECT 81.145 69.585 81.525 69.620 ;
        RECT 81.145 69.260 81.335 69.585 ;
        RECT 81.725 69.460 81.915 70.280 ;
        RECT 82.710 69.775 82.940 70.120 ;
        RECT 82.545 69.620 82.940 69.775 ;
        RECT 82.545 69.585 82.925 69.620 ;
        RECT 80.160 68.485 81.335 69.260 ;
        RECT 81.590 69.390 82.050 69.460 ;
        RECT 81.590 69.230 82.075 69.390 ;
        RECT 81.725 69.165 82.075 69.230 ;
        RECT 82.545 69.165 82.735 69.585 ;
        RECT 83.125 69.460 83.315 70.280 ;
        RECT 82.990 69.330 83.450 69.460 ;
        RECT 82.990 69.230 83.470 69.330 ;
        RECT 85.140 69.270 85.335 70.420 ;
        RECT 85.945 70.260 86.135 72.580 ;
        RECT 87.440 72.570 88.775 73.350 ;
        RECT 87.825 72.180 88.775 72.570 ;
        RECT 88.955 73.510 89.270 73.765 ;
        RECT 88.955 72.420 89.145 73.510 ;
        RECT 89.705 73.350 89.895 75.670 ;
        RECT 90.330 75.460 90.560 75.510 ;
        RECT 90.920 75.460 91.150 75.510 ;
        RECT 90.330 75.270 91.150 75.460 ;
        RECT 90.330 73.750 90.560 75.270 ;
        RECT 90.920 73.750 91.150 75.270 ;
        RECT 90.330 73.510 91.150 73.750 ;
        RECT 89.320 72.580 90.280 73.350 ;
        RECT 88.955 72.180 89.270 72.420 ;
        RECT 87.825 70.670 88.015 72.180 ;
        RECT 88.450 70.670 88.680 72.180 ;
        RECT 89.040 71.030 89.270 72.180 ;
        RECT 87.820 70.665 88.760 70.670 ;
        RECT 87.820 70.260 88.765 70.665 ;
        RECT 85.560 70.240 86.520 70.260 ;
        RECT 87.440 70.240 88.765 70.260 ;
        RECT 85.560 70.050 88.765 70.240 ;
        RECT 85.560 70.030 86.520 70.050 ;
        RECT 87.440 70.030 88.765 70.050 ;
        RECT 85.560 69.475 86.520 69.705 ;
        RECT 87.440 69.475 88.400 69.705 ;
        RECT 81.725 68.975 82.735 69.165 ;
        RECT 81.725 68.895 82.075 68.975 ;
        RECT 81.590 68.815 82.075 68.895 ;
        RECT 81.590 68.665 82.050 68.815 ;
        RECT 80.160 68.460 81.520 68.485 ;
        RECT 80.160 68.260 81.540 68.460 ;
        RECT 81.310 67.460 81.540 68.260 ;
        RECT 81.725 67.255 81.915 68.665 ;
        RECT 82.545 68.485 82.735 68.975 ;
        RECT 83.125 69.175 83.470 69.230 ;
        RECT 83.910 69.175 84.910 69.260 ;
        RECT 83.125 68.985 84.910 69.175 ;
        RECT 83.125 68.895 83.470 68.985 ;
        RECT 82.990 68.860 83.470 68.895 ;
        RECT 82.990 68.665 83.450 68.860 ;
        RECT 82.545 68.460 82.925 68.485 ;
        RECT 82.545 68.295 82.940 68.460 ;
        RECT 82.710 67.460 82.940 68.295 ;
        RECT 83.125 67.255 83.315 68.665 ;
        RECT 83.910 68.260 84.910 68.985 ;
        RECT 85.140 68.670 85.740 69.270 ;
        RECT 81.590 67.025 82.050 67.255 ;
        RECT 82.990 67.025 83.450 67.255 ;
        RECT 73.310 65.510 73.625 65.515 ;
        RECT 71.430 65.270 71.745 65.475 ;
        RECT 66.660 64.290 67.620 65.070 ;
        RECT 68.540 64.290 69.865 65.070 ;
        RECT 70.400 64.290 71.400 65.070 ;
        RECT 66.275 63.850 66.610 64.090 ;
        RECT 65.790 60.090 66.020 63.845 ;
        RECT 66.380 60.090 66.610 63.850 ;
        RECT 67.045 59.890 67.235 64.290 ;
        RECT 68.925 63.845 69.865 64.290 ;
        RECT 68.925 63.840 69.860 63.845 ;
        RECT 68.925 60.320 69.115 63.840 ;
        RECT 69.550 60.320 69.780 63.840 ;
        RECT 68.925 60.090 69.780 60.320 ;
        RECT 68.925 59.890 69.750 60.090 ;
        RECT 62.900 59.655 63.860 59.885 ;
        RECT 64.780 59.655 65.740 59.885 ;
        RECT 66.660 59.560 67.620 59.890 ;
        RECT 68.540 59.870 69.750 59.890 ;
        RECT 70.805 59.885 70.995 64.290 ;
        RECT 71.555 64.090 71.745 65.270 ;
        RECT 72.685 65.070 73.625 65.510 ;
        RECT 72.280 64.290 73.625 65.070 ;
        RECT 78.880 64.780 79.230 67.000 ;
        RECT 85.280 65.515 85.510 68.670 ;
        RECT 85.195 65.270 85.510 65.515 ;
        RECT 71.430 63.850 71.745 64.090 ;
        RECT 72.685 63.850 73.625 64.290 ;
        RECT 85.195 64.090 85.385 65.270 ;
        RECT 85.945 65.065 86.135 69.475 ;
        RECT 86.570 69.220 86.800 69.270 ;
        RECT 87.160 69.220 87.390 69.270 ;
        RECT 86.570 69.030 87.390 69.220 ;
        RECT 86.570 65.515 86.800 69.030 ;
        RECT 86.570 65.510 86.915 65.515 ;
        RECT 87.160 65.510 87.390 69.030 ;
        RECT 86.570 65.270 87.390 65.510 ;
        RECT 85.560 64.835 86.520 65.065 ;
        RECT 85.620 64.525 86.460 64.835 ;
        RECT 86.725 64.780 87.265 65.270 ;
        RECT 87.825 65.065 88.015 69.475 ;
        RECT 88.575 69.270 88.765 70.030 ;
        RECT 88.450 69.025 88.765 69.270 ;
        RECT 88.940 70.430 89.550 71.030 ;
        RECT 88.940 70.420 89.270 70.430 ;
        RECT 88.940 69.270 89.130 70.420 ;
        RECT 89.705 70.260 89.895 72.580 ;
        RECT 90.465 72.420 91.025 73.510 ;
        RECT 91.585 73.350 91.775 75.670 ;
        RECT 92.210 73.750 92.440 75.510 ;
        RECT 92.210 73.510 92.525 73.750 ;
        RECT 91.200 72.580 92.160 73.350 ;
        RECT 90.330 72.180 91.150 72.420 ;
        RECT 90.330 70.660 90.560 72.180 ;
        RECT 90.920 70.660 91.150 72.180 ;
        RECT 90.330 70.470 91.150 70.660 ;
        RECT 90.330 70.420 90.560 70.470 ;
        RECT 90.920 70.420 91.150 70.470 ;
        RECT 91.585 70.260 91.775 72.580 ;
        RECT 92.335 72.420 92.525 73.510 ;
        RECT 93.465 73.350 93.655 75.670 ;
        RECT 94.090 73.755 94.320 75.510 ;
        RECT 94.090 73.510 94.405 73.755 ;
        RECT 93.060 72.580 94.060 73.350 ;
        RECT 92.210 72.175 92.525 72.420 ;
        RECT 92.210 70.665 92.440 72.175 ;
        RECT 92.210 70.420 92.535 70.665 ;
        RECT 89.320 70.030 90.280 70.260 ;
        RECT 91.200 70.030 92.160 70.260 ;
        RECT 92.345 69.710 92.535 70.420 ;
        RECT 93.465 70.260 93.655 72.580 ;
        RECT 94.215 72.420 94.405 73.510 ;
        RECT 95.345 73.350 95.535 75.670 ;
        RECT 95.970 73.765 96.200 75.510 ;
        RECT 97.220 75.270 98.080 75.670 ;
        RECT 108.250 75.630 109.150 75.670 ;
        RECT 110.130 75.630 111.320 75.670 ;
        RECT 95.970 73.510 96.285 73.765 ;
        RECT 94.940 72.580 95.940 73.350 ;
        RECT 94.090 72.175 94.405 72.420 ;
        RECT 94.090 71.030 94.320 72.175 ;
        RECT 93.910 70.430 94.510 71.030 ;
        RECT 94.090 70.420 94.320 70.430 ;
        RECT 95.345 70.260 95.535 72.580 ;
        RECT 96.095 72.420 96.285 73.510 ;
        RECT 97.220 73.740 97.415 75.270 ;
        RECT 97.850 73.750 98.080 75.270 ;
        RECT 97.850 73.740 98.175 73.750 ;
        RECT 97.220 73.350 98.175 73.740 ;
        RECT 96.820 72.580 98.175 73.350 ;
        RECT 98.730 73.015 99.380 73.200 ;
        RECT 100.330 73.015 100.650 73.050 ;
        RECT 98.730 72.825 100.650 73.015 ;
        RECT 98.730 72.650 99.380 72.825 ;
        RECT 100.330 72.790 100.650 72.825 ;
        RECT 95.970 72.180 96.285 72.420 ;
        RECT 95.970 71.030 96.200 72.180 ;
        RECT 97.220 72.175 98.175 72.580 ;
        RECT 101.540 72.570 101.890 74.790 ;
        RECT 107.940 73.745 108.170 75.510 ;
        RECT 107.855 73.510 108.170 73.745 ;
        RECT 107.855 72.420 108.045 73.510 ;
        RECT 108.605 73.350 108.795 75.630 ;
        RECT 110.480 75.510 111.320 75.630 ;
        RECT 110.480 75.280 111.340 75.510 ;
        RECT 110.485 73.750 110.675 75.280 ;
        RECT 111.110 73.755 111.340 75.280 ;
        RECT 111.700 73.765 111.930 75.510 ;
        RECT 111.110 73.750 111.435 73.755 ;
        RECT 110.485 73.350 111.435 73.750 ;
        RECT 108.220 72.580 109.180 73.350 ;
        RECT 97.220 72.170 98.170 72.175 ;
        RECT 95.790 70.430 96.390 71.030 ;
        RECT 97.220 70.650 97.415 72.170 ;
        RECT 97.850 70.650 98.080 72.170 ;
        RECT 104.180 71.795 104.510 72.200 ;
        RECT 104.780 71.795 105.110 72.200 ;
        RECT 105.380 71.795 105.710 72.200 ;
        RECT 105.980 71.795 106.310 72.200 ;
        RECT 107.855 72.180 108.170 72.420 ;
        RECT 95.970 70.420 96.200 70.430 ;
        RECT 97.220 70.260 98.080 70.650 ;
        RECT 102.855 71.545 106.310 71.795 ;
        RECT 93.060 70.030 98.080 70.260 ;
        RECT 89.320 69.480 92.535 69.710 ;
        RECT 89.320 69.475 90.280 69.480 ;
        RECT 91.200 69.475 92.535 69.480 ;
        RECT 93.080 69.475 94.040 69.705 ;
        RECT 94.960 69.670 95.920 69.705 ;
        RECT 94.960 69.475 96.170 69.670 ;
        RECT 88.940 69.260 89.270 69.270 ;
        RECT 88.450 65.505 88.680 69.025 ;
        RECT 88.940 68.660 89.550 69.260 ;
        RECT 89.040 65.505 89.270 68.660 ;
        RECT 88.450 65.270 88.765 65.505 ;
        RECT 87.440 64.835 88.400 65.065 ;
        RECT 86.715 64.590 87.265 64.780 ;
        RECT 85.560 64.295 86.520 64.525 ;
        RECT 85.195 63.850 85.510 64.090 ;
        RECT 71.430 60.090 71.660 63.850 ;
        RECT 72.685 60.320 72.875 63.850 ;
        RECT 73.310 63.845 73.625 63.850 ;
        RECT 73.310 60.320 73.540 63.845 ;
        RECT 72.680 59.885 73.540 60.320 ;
        RECT 68.540 59.660 69.630 59.870 ;
        RECT 68.540 59.560 69.500 59.660 ;
        RECT 70.420 59.655 71.380 59.885 ;
        RECT 72.300 59.660 73.540 59.885 ;
        RECT 72.300 59.655 73.260 59.660 ;
        RECT 74.040 59.090 75.230 61.250 ;
        RECT 75.700 59.090 76.890 61.250 ;
        RECT 78.880 60.280 79.230 62.500 ;
        RECT 85.280 60.090 85.510 63.850 ;
        RECT 85.945 59.885 86.135 64.295 ;
        RECT 86.725 64.090 87.265 64.590 ;
        RECT 87.450 64.525 88.390 64.835 ;
        RECT 87.440 64.295 88.400 64.525 ;
        RECT 86.570 63.855 87.390 64.090 ;
        RECT 86.570 63.850 86.915 63.855 ;
        RECT 86.570 60.330 86.800 63.850 ;
        RECT 87.160 60.330 87.390 63.855 ;
        RECT 86.570 60.140 87.390 60.330 ;
        RECT 86.570 60.090 86.800 60.140 ;
        RECT 87.160 60.090 87.390 60.140 ;
        RECT 87.825 59.885 88.015 64.295 ;
        RECT 88.575 64.090 88.765 65.270 ;
        RECT 88.450 63.845 88.765 64.090 ;
        RECT 88.935 65.270 89.270 65.505 ;
        RECT 88.935 64.090 89.125 65.270 ;
        RECT 89.705 65.070 89.895 69.475 ;
        RECT 91.580 69.040 92.535 69.475 ;
        RECT 91.585 65.510 91.775 69.040 ;
        RECT 92.210 69.030 92.535 69.040 ;
        RECT 92.210 65.510 92.440 69.030 ;
        RECT 91.585 65.505 92.520 65.510 ;
        RECT 91.585 65.500 92.525 65.505 ;
        RECT 91.580 65.070 92.525 65.500 ;
        RECT 93.465 65.070 93.655 69.475 ;
        RECT 95.340 69.330 96.170 69.475 ;
        RECT 93.900 68.730 94.510 69.330 ;
        RECT 95.340 69.040 96.390 69.330 ;
        RECT 94.090 65.475 94.320 68.730 ;
        RECT 95.345 65.510 95.535 69.040 ;
        RECT 95.780 68.730 96.390 69.040 ;
        RECT 95.970 65.515 96.200 68.730 ;
        RECT 96.760 67.365 97.010 70.030 ;
        RECT 97.530 67.340 98.720 69.500 ;
        RECT 101.540 68.070 101.890 70.290 ;
        RECT 102.855 69.260 103.105 71.545 ;
        RECT 104.180 71.140 104.510 71.545 ;
        RECT 104.780 71.140 105.110 71.545 ;
        RECT 105.380 71.140 105.710 71.545 ;
        RECT 105.980 71.140 106.310 71.545 ;
        RECT 107.940 71.030 108.170 72.180 ;
        RECT 104.250 70.280 104.710 70.510 ;
        RECT 105.650 70.280 106.110 70.510 ;
        RECT 107.800 70.420 108.400 71.030 ;
        RECT 103.970 69.775 104.200 70.120 ;
        RECT 103.805 69.620 104.200 69.775 ;
        RECT 103.805 69.585 104.185 69.620 ;
        RECT 103.805 69.260 103.995 69.585 ;
        RECT 104.385 69.460 104.575 70.280 ;
        RECT 105.370 69.775 105.600 70.120 ;
        RECT 105.205 69.620 105.600 69.775 ;
        RECT 105.205 69.585 105.585 69.620 ;
        RECT 102.820 68.485 103.995 69.260 ;
        RECT 104.250 69.390 104.710 69.460 ;
        RECT 104.250 69.230 104.735 69.390 ;
        RECT 104.385 69.165 104.735 69.230 ;
        RECT 105.205 69.165 105.395 69.585 ;
        RECT 105.785 69.460 105.975 70.280 ;
        RECT 105.650 69.330 106.110 69.460 ;
        RECT 105.650 69.230 106.130 69.330 ;
        RECT 107.800 69.270 107.995 70.420 ;
        RECT 108.605 70.260 108.795 72.580 ;
        RECT 110.100 72.570 111.435 73.350 ;
        RECT 110.485 72.180 111.435 72.570 ;
        RECT 111.615 73.510 111.930 73.765 ;
        RECT 111.615 72.420 111.805 73.510 ;
        RECT 112.365 73.350 112.555 75.670 ;
        RECT 112.990 75.460 113.220 75.510 ;
        RECT 113.580 75.460 113.810 75.510 ;
        RECT 112.990 75.270 113.810 75.460 ;
        RECT 112.990 73.750 113.220 75.270 ;
        RECT 113.580 73.750 113.810 75.270 ;
        RECT 112.990 73.510 113.810 73.750 ;
        RECT 111.980 72.580 112.940 73.350 ;
        RECT 111.615 72.180 111.930 72.420 ;
        RECT 110.485 70.670 110.675 72.180 ;
        RECT 111.110 70.670 111.340 72.180 ;
        RECT 111.700 71.030 111.930 72.180 ;
        RECT 110.480 70.665 111.420 70.670 ;
        RECT 110.480 70.260 111.425 70.665 ;
        RECT 108.220 70.240 109.180 70.260 ;
        RECT 110.100 70.240 111.425 70.260 ;
        RECT 108.220 70.050 111.425 70.240 ;
        RECT 108.220 70.030 109.180 70.050 ;
        RECT 110.100 70.030 111.425 70.050 ;
        RECT 108.220 69.475 109.180 69.705 ;
        RECT 110.100 69.475 111.060 69.705 ;
        RECT 104.385 68.975 105.395 69.165 ;
        RECT 104.385 68.895 104.735 68.975 ;
        RECT 104.250 68.815 104.735 68.895 ;
        RECT 104.250 68.665 104.710 68.815 ;
        RECT 102.820 68.460 104.180 68.485 ;
        RECT 102.820 68.260 104.200 68.460 ;
        RECT 103.970 67.460 104.200 68.260 ;
        RECT 104.385 67.255 104.575 68.665 ;
        RECT 105.205 68.485 105.395 68.975 ;
        RECT 105.785 69.175 106.130 69.230 ;
        RECT 106.570 69.175 107.570 69.260 ;
        RECT 105.785 68.985 107.570 69.175 ;
        RECT 105.785 68.895 106.130 68.985 ;
        RECT 105.650 68.860 106.130 68.895 ;
        RECT 105.650 68.665 106.110 68.860 ;
        RECT 105.205 68.460 105.585 68.485 ;
        RECT 105.205 68.295 105.600 68.460 ;
        RECT 105.370 67.460 105.600 68.295 ;
        RECT 105.785 67.255 105.975 68.665 ;
        RECT 106.570 68.260 107.570 68.985 ;
        RECT 107.800 68.670 108.400 69.270 ;
        RECT 104.250 67.025 104.710 67.255 ;
        RECT 105.650 67.025 106.110 67.255 ;
        RECT 95.970 65.510 96.285 65.515 ;
        RECT 94.090 65.270 94.405 65.475 ;
        RECT 89.320 64.290 90.280 65.070 ;
        RECT 91.200 64.290 92.525 65.070 ;
        RECT 93.060 64.290 94.060 65.070 ;
        RECT 88.935 63.850 89.270 64.090 ;
        RECT 88.450 60.090 88.680 63.845 ;
        RECT 89.040 60.090 89.270 63.850 ;
        RECT 89.705 59.890 89.895 64.290 ;
        RECT 91.585 63.845 92.525 64.290 ;
        RECT 91.585 63.840 92.520 63.845 ;
        RECT 91.585 60.320 91.775 63.840 ;
        RECT 92.210 60.320 92.440 63.840 ;
        RECT 91.585 60.090 92.440 60.320 ;
        RECT 91.585 59.890 92.410 60.090 ;
        RECT 85.560 59.655 86.520 59.885 ;
        RECT 87.440 59.655 88.400 59.885 ;
        RECT 89.320 59.560 90.280 59.890 ;
        RECT 91.200 59.870 92.410 59.890 ;
        RECT 93.465 59.885 93.655 64.290 ;
        RECT 94.215 64.090 94.405 65.270 ;
        RECT 95.345 65.070 96.285 65.510 ;
        RECT 94.940 64.290 96.285 65.070 ;
        RECT 101.540 64.780 101.890 67.000 ;
        RECT 107.940 65.515 108.170 68.670 ;
        RECT 107.855 65.270 108.170 65.515 ;
        RECT 94.090 63.850 94.405 64.090 ;
        RECT 95.345 63.850 96.285 64.290 ;
        RECT 107.855 64.090 108.045 65.270 ;
        RECT 108.605 65.065 108.795 69.475 ;
        RECT 109.230 69.220 109.460 69.270 ;
        RECT 109.820 69.220 110.050 69.270 ;
        RECT 109.230 69.030 110.050 69.220 ;
        RECT 109.230 65.515 109.460 69.030 ;
        RECT 109.230 65.510 109.575 65.515 ;
        RECT 109.820 65.510 110.050 69.030 ;
        RECT 109.230 65.270 110.050 65.510 ;
        RECT 108.220 64.835 109.180 65.065 ;
        RECT 108.280 64.525 109.120 64.835 ;
        RECT 109.385 64.780 109.925 65.270 ;
        RECT 110.485 65.065 110.675 69.475 ;
        RECT 111.235 69.270 111.425 70.030 ;
        RECT 111.110 69.025 111.425 69.270 ;
        RECT 111.600 70.430 112.210 71.030 ;
        RECT 111.600 70.420 111.930 70.430 ;
        RECT 111.600 69.270 111.790 70.420 ;
        RECT 112.365 70.260 112.555 72.580 ;
        RECT 113.125 72.420 113.685 73.510 ;
        RECT 114.245 73.350 114.435 75.670 ;
        RECT 114.870 73.750 115.100 75.510 ;
        RECT 114.870 73.510 115.185 73.750 ;
        RECT 113.860 72.580 114.820 73.350 ;
        RECT 112.990 72.180 113.810 72.420 ;
        RECT 112.990 70.660 113.220 72.180 ;
        RECT 113.580 70.660 113.810 72.180 ;
        RECT 112.990 70.470 113.810 70.660 ;
        RECT 112.990 70.420 113.220 70.470 ;
        RECT 113.580 70.420 113.810 70.470 ;
        RECT 114.245 70.260 114.435 72.580 ;
        RECT 114.995 72.420 115.185 73.510 ;
        RECT 116.125 73.350 116.315 75.670 ;
        RECT 116.750 73.755 116.980 75.510 ;
        RECT 116.750 73.510 117.065 73.755 ;
        RECT 115.720 72.580 116.720 73.350 ;
        RECT 114.870 72.175 115.185 72.420 ;
        RECT 114.870 70.665 115.100 72.175 ;
        RECT 114.870 70.420 115.195 70.665 ;
        RECT 111.980 70.030 112.940 70.260 ;
        RECT 113.860 70.030 114.820 70.260 ;
        RECT 115.005 69.710 115.195 70.420 ;
        RECT 116.125 70.260 116.315 72.580 ;
        RECT 116.875 72.420 117.065 73.510 ;
        RECT 118.005 73.350 118.195 75.670 ;
        RECT 118.630 73.765 118.860 75.510 ;
        RECT 119.880 75.270 120.740 75.670 ;
        RECT 118.630 73.510 118.945 73.765 ;
        RECT 117.600 72.580 118.600 73.350 ;
        RECT 116.750 72.175 117.065 72.420 ;
        RECT 116.750 71.030 116.980 72.175 ;
        RECT 116.570 70.430 117.170 71.030 ;
        RECT 116.750 70.420 116.980 70.430 ;
        RECT 118.005 70.260 118.195 72.580 ;
        RECT 118.755 72.420 118.945 73.510 ;
        RECT 119.880 73.740 120.075 75.270 ;
        RECT 120.510 73.750 120.740 75.270 ;
        RECT 120.510 73.740 120.835 73.750 ;
        RECT 119.880 73.350 120.835 73.740 ;
        RECT 119.480 72.580 120.835 73.350 ;
        RECT 121.390 73.015 122.040 73.200 ;
        RECT 122.990 73.015 123.310 73.050 ;
        RECT 121.390 72.825 123.310 73.015 ;
        RECT 121.390 72.650 122.040 72.825 ;
        RECT 122.990 72.790 123.310 72.825 ;
        RECT 118.630 72.180 118.945 72.420 ;
        RECT 118.630 71.030 118.860 72.180 ;
        RECT 119.880 72.175 120.835 72.580 ;
        RECT 124.200 72.570 124.550 74.790 ;
        RECT 119.880 72.170 120.830 72.175 ;
        RECT 118.450 70.430 119.050 71.030 ;
        RECT 119.880 70.650 120.075 72.170 ;
        RECT 120.510 70.650 120.740 72.170 ;
        RECT 118.630 70.420 118.860 70.430 ;
        RECT 119.880 70.260 120.740 70.650 ;
        RECT 115.720 70.030 120.740 70.260 ;
        RECT 111.980 69.480 115.195 69.710 ;
        RECT 111.980 69.475 112.940 69.480 ;
        RECT 113.860 69.475 115.195 69.480 ;
        RECT 115.740 69.475 116.700 69.705 ;
        RECT 117.620 69.670 118.580 69.705 ;
        RECT 117.620 69.475 118.830 69.670 ;
        RECT 111.600 69.260 111.930 69.270 ;
        RECT 111.110 65.505 111.340 69.025 ;
        RECT 111.600 68.660 112.210 69.260 ;
        RECT 111.700 65.505 111.930 68.660 ;
        RECT 111.110 65.270 111.425 65.505 ;
        RECT 110.100 64.835 111.060 65.065 ;
        RECT 109.375 64.590 109.925 64.780 ;
        RECT 108.220 64.295 109.180 64.525 ;
        RECT 107.855 63.850 108.170 64.090 ;
        RECT 94.090 60.090 94.320 63.850 ;
        RECT 95.345 60.320 95.535 63.850 ;
        RECT 95.970 63.845 96.285 63.850 ;
        RECT 95.970 60.320 96.200 63.845 ;
        RECT 95.340 59.885 96.200 60.320 ;
        RECT 91.200 59.660 92.290 59.870 ;
        RECT 91.200 59.560 92.160 59.660 ;
        RECT 93.080 59.655 94.040 59.885 ;
        RECT 94.960 59.660 96.200 59.885 ;
        RECT 94.960 59.655 95.920 59.660 ;
        RECT 96.700 59.090 97.890 61.250 ;
        RECT 98.360 59.090 99.550 61.250 ;
        RECT 101.540 60.280 101.890 62.500 ;
        RECT 107.940 60.090 108.170 63.850 ;
        RECT 108.605 59.885 108.795 64.295 ;
        RECT 109.385 64.090 109.925 64.590 ;
        RECT 110.110 64.525 111.050 64.835 ;
        RECT 110.100 64.295 111.060 64.525 ;
        RECT 109.230 63.855 110.050 64.090 ;
        RECT 109.230 63.850 109.575 63.855 ;
        RECT 109.230 60.330 109.460 63.850 ;
        RECT 109.820 60.330 110.050 63.855 ;
        RECT 109.230 60.140 110.050 60.330 ;
        RECT 109.230 60.090 109.460 60.140 ;
        RECT 109.820 60.090 110.050 60.140 ;
        RECT 110.485 59.885 110.675 64.295 ;
        RECT 111.235 64.090 111.425 65.270 ;
        RECT 111.110 63.845 111.425 64.090 ;
        RECT 111.595 65.270 111.930 65.505 ;
        RECT 111.595 64.090 111.785 65.270 ;
        RECT 112.365 65.070 112.555 69.475 ;
        RECT 114.240 69.040 115.195 69.475 ;
        RECT 114.245 65.510 114.435 69.040 ;
        RECT 114.870 69.030 115.195 69.040 ;
        RECT 114.870 65.510 115.100 69.030 ;
        RECT 114.245 65.505 115.180 65.510 ;
        RECT 114.245 65.500 115.185 65.505 ;
        RECT 114.240 65.070 115.185 65.500 ;
        RECT 116.125 65.070 116.315 69.475 ;
        RECT 118.000 69.330 118.830 69.475 ;
        RECT 116.560 68.730 117.170 69.330 ;
        RECT 118.000 69.040 119.050 69.330 ;
        RECT 116.750 65.475 116.980 68.730 ;
        RECT 118.005 65.510 118.195 69.040 ;
        RECT 118.440 68.730 119.050 69.040 ;
        RECT 118.630 65.515 118.860 68.730 ;
        RECT 119.420 67.365 119.670 70.030 ;
        RECT 120.190 67.340 121.380 69.500 ;
        RECT 124.200 68.070 124.550 70.290 ;
        RECT 118.630 65.510 118.945 65.515 ;
        RECT 116.750 65.270 117.065 65.475 ;
        RECT 111.980 64.290 112.940 65.070 ;
        RECT 113.860 64.290 115.185 65.070 ;
        RECT 115.720 64.290 116.720 65.070 ;
        RECT 111.595 63.850 111.930 64.090 ;
        RECT 111.110 60.090 111.340 63.845 ;
        RECT 111.700 60.090 111.930 63.850 ;
        RECT 112.365 59.890 112.555 64.290 ;
        RECT 114.245 63.845 115.185 64.290 ;
        RECT 114.245 63.840 115.180 63.845 ;
        RECT 114.245 60.320 114.435 63.840 ;
        RECT 114.870 60.320 115.100 63.840 ;
        RECT 114.245 60.090 115.100 60.320 ;
        RECT 114.245 59.890 115.070 60.090 ;
        RECT 108.220 59.655 109.180 59.885 ;
        RECT 110.100 59.655 111.060 59.885 ;
        RECT 111.980 59.560 112.940 59.890 ;
        RECT 113.860 59.870 115.070 59.890 ;
        RECT 116.125 59.885 116.315 64.290 ;
        RECT 116.875 64.090 117.065 65.270 ;
        RECT 118.005 65.070 118.945 65.510 ;
        RECT 117.600 64.290 118.945 65.070 ;
        RECT 124.200 64.780 124.550 67.000 ;
        RECT 116.750 63.850 117.065 64.090 ;
        RECT 118.005 63.850 118.945 64.290 ;
        RECT 116.750 60.090 116.980 63.850 ;
        RECT 118.005 60.320 118.195 63.850 ;
        RECT 118.630 63.845 118.945 63.850 ;
        RECT 118.630 60.320 118.860 63.845 ;
        RECT 118.000 59.885 118.860 60.320 ;
        RECT 113.860 59.660 114.950 59.870 ;
        RECT 113.860 59.560 114.820 59.660 ;
        RECT 115.740 59.655 116.700 59.885 ;
        RECT 117.620 59.660 118.860 59.885 ;
        RECT 117.620 59.655 118.580 59.660 ;
        RECT 119.360 59.090 120.550 61.250 ;
        RECT 121.020 59.090 122.210 61.250 ;
        RECT 124.200 60.280 124.550 62.500 ;
        RECT 56.230 58.875 56.550 58.880 ;
        RECT 78.900 58.875 79.220 58.880 ;
        RECT 56.230 58.625 79.220 58.875 ;
        RECT 56.230 58.620 56.550 58.625 ;
        RECT 78.900 58.620 79.220 58.625 ;
        RECT 101.555 58.875 101.875 58.880 ;
        RECT 124.215 58.875 124.535 58.880 ;
        RECT 101.555 58.625 124.535 58.875 ;
        RECT 101.555 58.620 101.875 58.625 ;
        RECT 124.215 58.620 124.535 58.625 ;
        RECT 40.270 57.900 41.170 57.950 ;
        RECT 42.150 57.900 43.050 57.950 ;
        RECT 40.240 57.670 41.200 57.900 ;
        RECT 42.120 57.875 43.080 57.900 ;
        RECT 42.120 57.670 43.340 57.875 ;
        RECT 44.000 57.670 44.960 57.900 ;
        RECT 47.740 57.670 48.740 57.990 ;
        RECT 49.620 57.670 50.620 57.990 ;
        RECT 51.500 57.900 52.500 57.990 ;
        RECT 62.930 57.900 63.830 57.950 ;
        RECT 64.810 57.900 65.710 57.950 ;
        RECT 51.500 57.670 52.760 57.900 ;
        RECT 62.900 57.670 63.860 57.900 ;
        RECT 64.780 57.875 65.740 57.900 ;
        RECT 64.780 57.670 66.000 57.875 ;
        RECT 66.660 57.670 67.620 57.900 ;
        RECT 70.400 57.670 71.400 57.990 ;
        RECT 72.280 57.670 73.280 57.990 ;
        RECT 74.160 57.900 75.160 57.990 ;
        RECT 85.590 57.900 86.490 57.950 ;
        RECT 87.470 57.900 88.370 57.950 ;
        RECT 74.160 57.670 75.420 57.900 ;
        RECT 85.560 57.670 86.520 57.900 ;
        RECT 87.440 57.875 88.400 57.900 ;
        RECT 87.440 57.670 88.660 57.875 ;
        RECT 89.320 57.670 90.280 57.900 ;
        RECT 93.060 57.670 94.060 57.990 ;
        RECT 94.940 57.670 95.940 57.990 ;
        RECT 96.820 57.900 97.820 57.990 ;
        RECT 108.250 57.900 109.150 57.950 ;
        RECT 110.130 57.900 111.030 57.950 ;
        RECT 96.820 57.670 98.080 57.900 ;
        RECT 108.220 57.670 109.180 57.900 ;
        RECT 110.100 57.875 111.060 57.900 ;
        RECT 110.100 57.670 111.320 57.875 ;
        RECT 111.980 57.670 112.940 57.900 ;
        RECT 115.720 57.670 116.720 57.990 ;
        RECT 117.600 57.670 118.600 57.990 ;
        RECT 119.480 57.900 120.480 57.990 ;
        RECT 119.480 57.670 120.740 57.900 ;
        RECT 40.270 57.630 41.170 57.670 ;
        RECT 42.150 57.630 43.340 57.670 ;
        RECT 39.960 55.745 40.190 57.510 ;
        RECT 39.875 55.510 40.190 55.745 ;
        RECT 39.875 54.420 40.065 55.510 ;
        RECT 40.625 55.350 40.815 57.630 ;
        RECT 42.500 57.510 43.340 57.630 ;
        RECT 42.500 57.280 43.360 57.510 ;
        RECT 42.505 55.750 42.695 57.280 ;
        RECT 43.130 55.755 43.360 57.280 ;
        RECT 43.720 55.765 43.950 57.510 ;
        RECT 43.130 55.750 43.455 55.755 ;
        RECT 42.505 55.350 43.455 55.750 ;
        RECT 40.240 54.580 41.200 55.350 ;
        RECT 39.875 54.180 40.190 54.420 ;
        RECT 39.960 53.030 40.190 54.180 ;
        RECT 39.820 52.420 40.420 53.030 ;
        RECT 39.820 51.270 40.015 52.420 ;
        RECT 40.625 52.260 40.815 54.580 ;
        RECT 42.120 54.570 43.455 55.350 ;
        RECT 42.505 54.180 43.455 54.570 ;
        RECT 43.635 55.510 43.950 55.765 ;
        RECT 43.635 54.420 43.825 55.510 ;
        RECT 44.385 55.350 44.575 57.670 ;
        RECT 45.010 57.460 45.240 57.510 ;
        RECT 45.600 57.460 45.830 57.510 ;
        RECT 45.010 57.270 45.830 57.460 ;
        RECT 45.010 55.750 45.240 57.270 ;
        RECT 45.600 55.750 45.830 57.270 ;
        RECT 45.010 55.510 45.830 55.750 ;
        RECT 46.890 55.750 47.120 57.510 ;
        RECT 46.890 55.510 47.205 55.750 ;
        RECT 44.000 54.580 44.960 55.350 ;
        RECT 43.635 54.180 43.950 54.420 ;
        RECT 42.505 52.670 42.695 54.180 ;
        RECT 43.130 52.670 43.360 54.180 ;
        RECT 43.720 53.030 43.950 54.180 ;
        RECT 42.500 52.665 43.440 52.670 ;
        RECT 42.500 52.260 43.445 52.665 ;
        RECT 40.240 52.240 41.200 52.260 ;
        RECT 42.120 52.240 43.445 52.260 ;
        RECT 40.240 52.050 43.445 52.240 ;
        RECT 40.240 52.030 41.200 52.050 ;
        RECT 42.120 52.030 43.445 52.050 ;
        RECT 40.240 51.475 41.200 51.705 ;
        RECT 39.820 50.670 40.420 51.270 ;
        RECT 39.960 47.515 40.190 50.670 ;
        RECT 39.875 47.270 40.190 47.515 ;
        RECT 39.875 46.090 40.065 47.270 ;
        RECT 40.625 47.065 40.815 51.475 ;
        RECT 43.255 51.270 43.445 52.030 ;
        RECT 41.250 51.220 41.480 51.270 ;
        RECT 41.840 51.220 42.070 51.270 ;
        RECT 41.250 51.030 42.070 51.220 ;
        RECT 41.250 47.515 41.480 51.030 ;
        RECT 41.250 47.510 41.595 47.515 ;
        RECT 41.840 47.510 42.070 51.030 ;
        RECT 41.250 47.270 42.070 47.510 ;
        RECT 43.130 51.025 43.445 51.270 ;
        RECT 43.620 52.430 44.230 53.030 ;
        RECT 43.620 52.420 43.950 52.430 ;
        RECT 43.620 51.270 43.810 52.420 ;
        RECT 44.385 52.260 44.575 54.580 ;
        RECT 45.145 54.420 45.705 55.510 ;
        RECT 47.015 54.420 47.205 55.510 ;
        RECT 48.145 55.350 48.335 57.670 ;
        RECT 48.770 55.755 49.000 57.510 ;
        RECT 48.770 55.510 49.085 55.755 ;
        RECT 47.740 54.580 48.740 55.350 ;
        RECT 45.010 54.180 45.830 54.420 ;
        RECT 45.010 52.660 45.240 54.180 ;
        RECT 45.600 52.660 45.830 54.180 ;
        RECT 45.010 52.470 45.830 52.660 ;
        RECT 45.010 52.420 45.240 52.470 ;
        RECT 45.600 52.420 45.830 52.470 ;
        RECT 46.890 54.175 47.205 54.420 ;
        RECT 46.890 52.665 47.120 54.175 ;
        RECT 46.890 52.420 47.215 52.665 ;
        RECT 44.000 52.030 44.960 52.260 ;
        RECT 47.025 51.710 47.215 52.420 ;
        RECT 48.145 52.260 48.335 54.580 ;
        RECT 48.895 54.420 49.085 55.510 ;
        RECT 50.025 55.350 50.215 57.670 ;
        RECT 50.650 55.765 50.880 57.510 ;
        RECT 51.900 57.270 52.760 57.670 ;
        RECT 62.930 57.630 63.830 57.670 ;
        RECT 64.810 57.630 66.000 57.670 ;
        RECT 50.650 55.510 50.965 55.765 ;
        RECT 49.620 54.580 50.620 55.350 ;
        RECT 48.770 54.175 49.085 54.420 ;
        RECT 48.770 53.030 49.000 54.175 ;
        RECT 48.590 52.430 49.190 53.030 ;
        RECT 48.770 52.420 49.000 52.430 ;
        RECT 50.025 52.260 50.215 54.580 ;
        RECT 50.775 54.420 50.965 55.510 ;
        RECT 51.900 55.740 52.095 57.270 ;
        RECT 52.530 55.750 52.760 57.270 ;
        RECT 52.530 55.740 52.855 55.750 ;
        RECT 62.620 55.745 62.850 57.510 ;
        RECT 51.900 55.350 52.855 55.740 ;
        RECT 51.500 54.580 52.855 55.350 ;
        RECT 50.650 54.180 50.965 54.420 ;
        RECT 50.650 53.030 50.880 54.180 ;
        RECT 51.900 54.175 52.855 54.580 ;
        RECT 62.535 55.510 62.850 55.745 ;
        RECT 62.535 54.420 62.725 55.510 ;
        RECT 63.285 55.350 63.475 57.630 ;
        RECT 65.160 57.510 66.000 57.630 ;
        RECT 65.160 57.280 66.020 57.510 ;
        RECT 65.165 55.750 65.355 57.280 ;
        RECT 65.790 55.755 66.020 57.280 ;
        RECT 66.380 55.765 66.610 57.510 ;
        RECT 65.790 55.750 66.115 55.755 ;
        RECT 65.165 55.350 66.115 55.750 ;
        RECT 62.900 54.580 63.860 55.350 ;
        RECT 62.535 54.180 62.850 54.420 ;
        RECT 51.900 54.170 52.850 54.175 ;
        RECT 50.470 52.430 51.070 53.030 ;
        RECT 51.900 52.650 52.095 54.170 ;
        RECT 52.530 52.650 52.760 54.170 ;
        RECT 62.620 53.030 62.850 54.180 ;
        RECT 50.650 52.420 50.880 52.430 ;
        RECT 51.900 52.260 52.760 52.650 ;
        RECT 47.740 52.030 52.760 52.260 ;
        RECT 62.480 52.420 63.080 53.030 ;
        RECT 44.000 51.480 47.215 51.710 ;
        RECT 44.000 51.475 44.960 51.480 ;
        RECT 45.880 51.475 47.215 51.480 ;
        RECT 47.760 51.475 48.720 51.705 ;
        RECT 49.640 51.670 50.600 51.705 ;
        RECT 49.640 51.475 50.850 51.670 ;
        RECT 43.620 51.260 43.950 51.270 ;
        RECT 43.130 47.505 43.360 51.025 ;
        RECT 43.620 50.660 44.230 51.260 ;
        RECT 43.720 47.505 43.950 50.660 ;
        RECT 43.130 47.270 43.445 47.505 ;
        RECT 40.240 46.835 41.200 47.065 ;
        RECT 40.300 46.525 41.140 46.835 ;
        RECT 41.405 46.780 41.945 47.270 ;
        RECT 41.395 46.590 41.945 46.780 ;
        RECT 40.240 46.295 41.200 46.525 ;
        RECT 39.875 45.850 40.190 46.090 ;
        RECT 39.960 42.090 40.190 45.850 ;
        RECT 40.625 41.885 40.815 46.295 ;
        RECT 41.405 46.090 41.945 46.590 ;
        RECT 43.255 46.090 43.445 47.270 ;
        RECT 41.250 45.855 42.070 46.090 ;
        RECT 41.250 45.850 41.595 45.855 ;
        RECT 41.250 42.330 41.480 45.850 ;
        RECT 41.840 42.330 42.070 45.855 ;
        RECT 41.250 42.140 42.070 42.330 ;
        RECT 41.250 42.090 41.480 42.140 ;
        RECT 41.840 42.090 42.070 42.140 ;
        RECT 43.130 45.845 43.445 46.090 ;
        RECT 43.615 47.270 43.950 47.505 ;
        RECT 43.615 46.090 43.805 47.270 ;
        RECT 44.385 47.070 44.575 51.475 ;
        RECT 46.260 51.040 47.215 51.475 ;
        RECT 46.265 47.510 46.455 51.040 ;
        RECT 46.890 51.030 47.215 51.040 ;
        RECT 46.890 47.510 47.120 51.030 ;
        RECT 46.265 47.505 47.200 47.510 ;
        RECT 46.265 47.500 47.205 47.505 ;
        RECT 46.260 47.070 47.205 47.500 ;
        RECT 48.145 47.070 48.335 51.475 ;
        RECT 50.020 51.330 50.850 51.475 ;
        RECT 48.580 50.730 49.190 51.330 ;
        RECT 50.020 51.040 51.070 51.330 ;
        RECT 48.770 47.475 49.000 50.730 ;
        RECT 50.025 47.510 50.215 51.040 ;
        RECT 50.460 50.730 51.070 51.040 ;
        RECT 50.650 47.515 50.880 50.730 ;
        RECT 51.440 49.365 51.690 52.030 ;
        RECT 52.210 49.340 53.400 51.500 ;
        RECT 62.480 51.270 62.675 52.420 ;
        RECT 63.285 52.260 63.475 54.580 ;
        RECT 64.780 54.570 66.115 55.350 ;
        RECT 65.165 54.180 66.115 54.570 ;
        RECT 66.295 55.510 66.610 55.765 ;
        RECT 66.295 54.420 66.485 55.510 ;
        RECT 67.045 55.350 67.235 57.670 ;
        RECT 67.670 57.460 67.900 57.510 ;
        RECT 68.260 57.460 68.490 57.510 ;
        RECT 67.670 57.270 68.490 57.460 ;
        RECT 67.670 55.750 67.900 57.270 ;
        RECT 68.260 55.750 68.490 57.270 ;
        RECT 67.670 55.510 68.490 55.750 ;
        RECT 69.550 55.750 69.780 57.510 ;
        RECT 69.550 55.510 69.865 55.750 ;
        RECT 66.660 54.580 67.620 55.350 ;
        RECT 66.295 54.180 66.610 54.420 ;
        RECT 65.165 52.670 65.355 54.180 ;
        RECT 65.790 52.670 66.020 54.180 ;
        RECT 66.380 53.030 66.610 54.180 ;
        RECT 65.160 52.665 66.100 52.670 ;
        RECT 65.160 52.260 66.105 52.665 ;
        RECT 62.900 52.240 63.860 52.260 ;
        RECT 64.780 52.240 66.105 52.260 ;
        RECT 62.900 52.050 66.105 52.240 ;
        RECT 62.900 52.030 63.860 52.050 ;
        RECT 64.780 52.030 66.105 52.050 ;
        RECT 62.900 51.475 63.860 51.705 ;
        RECT 62.480 50.670 63.080 51.270 ;
        RECT 62.620 47.515 62.850 50.670 ;
        RECT 50.650 47.510 50.965 47.515 ;
        RECT 48.770 47.270 49.085 47.475 ;
        RECT 44.000 46.290 44.960 47.070 ;
        RECT 45.880 46.290 47.205 47.070 ;
        RECT 47.740 46.290 48.740 47.070 ;
        RECT 43.615 45.850 43.950 46.090 ;
        RECT 43.130 42.090 43.360 45.845 ;
        RECT 43.720 42.090 43.950 45.850 ;
        RECT 44.385 41.890 44.575 46.290 ;
        RECT 46.265 45.845 47.205 46.290 ;
        RECT 46.265 45.840 47.200 45.845 ;
        RECT 46.265 42.320 46.455 45.840 ;
        RECT 46.890 42.320 47.120 45.840 ;
        RECT 46.265 42.090 47.120 42.320 ;
        RECT 46.265 41.890 47.090 42.090 ;
        RECT 40.240 41.655 41.200 41.885 ;
        RECT 44.000 41.560 44.960 41.890 ;
        RECT 45.880 41.870 47.090 41.890 ;
        RECT 48.145 41.885 48.335 46.290 ;
        RECT 48.895 46.090 49.085 47.270 ;
        RECT 50.025 47.070 50.965 47.510 ;
        RECT 49.620 46.290 50.965 47.070 ;
        RECT 48.770 45.850 49.085 46.090 ;
        RECT 50.025 45.850 50.965 46.290 ;
        RECT 62.535 47.270 62.850 47.515 ;
        RECT 62.535 46.090 62.725 47.270 ;
        RECT 63.285 47.065 63.475 51.475 ;
        RECT 65.915 51.270 66.105 52.030 ;
        RECT 63.910 51.220 64.140 51.270 ;
        RECT 64.500 51.220 64.730 51.270 ;
        RECT 63.910 51.030 64.730 51.220 ;
        RECT 63.910 47.515 64.140 51.030 ;
        RECT 63.910 47.510 64.255 47.515 ;
        RECT 64.500 47.510 64.730 51.030 ;
        RECT 63.910 47.270 64.730 47.510 ;
        RECT 65.790 51.025 66.105 51.270 ;
        RECT 66.280 52.430 66.890 53.030 ;
        RECT 66.280 52.420 66.610 52.430 ;
        RECT 66.280 51.270 66.470 52.420 ;
        RECT 67.045 52.260 67.235 54.580 ;
        RECT 67.805 54.420 68.365 55.510 ;
        RECT 69.675 54.420 69.865 55.510 ;
        RECT 70.805 55.350 70.995 57.670 ;
        RECT 71.430 55.755 71.660 57.510 ;
        RECT 71.430 55.510 71.745 55.755 ;
        RECT 70.400 54.580 71.400 55.350 ;
        RECT 67.670 54.180 68.490 54.420 ;
        RECT 67.670 52.660 67.900 54.180 ;
        RECT 68.260 52.660 68.490 54.180 ;
        RECT 67.670 52.470 68.490 52.660 ;
        RECT 67.670 52.420 67.900 52.470 ;
        RECT 68.260 52.420 68.490 52.470 ;
        RECT 69.550 54.175 69.865 54.420 ;
        RECT 69.550 52.665 69.780 54.175 ;
        RECT 69.550 52.420 69.875 52.665 ;
        RECT 66.660 52.030 67.620 52.260 ;
        RECT 69.685 51.710 69.875 52.420 ;
        RECT 70.805 52.260 70.995 54.580 ;
        RECT 71.555 54.420 71.745 55.510 ;
        RECT 72.685 55.350 72.875 57.670 ;
        RECT 73.310 55.765 73.540 57.510 ;
        RECT 74.560 57.270 75.420 57.670 ;
        RECT 85.590 57.630 86.490 57.670 ;
        RECT 87.470 57.630 88.660 57.670 ;
        RECT 73.310 55.510 73.625 55.765 ;
        RECT 72.280 54.580 73.280 55.350 ;
        RECT 71.430 54.175 71.745 54.420 ;
        RECT 71.430 53.030 71.660 54.175 ;
        RECT 71.250 52.430 71.850 53.030 ;
        RECT 71.430 52.420 71.660 52.430 ;
        RECT 72.685 52.260 72.875 54.580 ;
        RECT 73.435 54.420 73.625 55.510 ;
        RECT 74.560 55.740 74.755 57.270 ;
        RECT 75.190 55.750 75.420 57.270 ;
        RECT 75.190 55.740 75.515 55.750 ;
        RECT 85.280 55.745 85.510 57.510 ;
        RECT 74.560 55.350 75.515 55.740 ;
        RECT 74.160 54.580 75.515 55.350 ;
        RECT 73.310 54.180 73.625 54.420 ;
        RECT 73.310 53.030 73.540 54.180 ;
        RECT 74.560 54.175 75.515 54.580 ;
        RECT 85.195 55.510 85.510 55.745 ;
        RECT 85.195 54.420 85.385 55.510 ;
        RECT 85.945 55.350 86.135 57.630 ;
        RECT 87.820 57.510 88.660 57.630 ;
        RECT 87.820 57.280 88.680 57.510 ;
        RECT 87.825 55.750 88.015 57.280 ;
        RECT 88.450 55.755 88.680 57.280 ;
        RECT 89.040 55.765 89.270 57.510 ;
        RECT 88.450 55.750 88.775 55.755 ;
        RECT 87.825 55.350 88.775 55.750 ;
        RECT 85.560 54.580 86.520 55.350 ;
        RECT 85.195 54.180 85.510 54.420 ;
        RECT 74.560 54.170 75.510 54.175 ;
        RECT 73.130 52.430 73.730 53.030 ;
        RECT 74.560 52.650 74.755 54.170 ;
        RECT 75.190 52.650 75.420 54.170 ;
        RECT 85.280 53.030 85.510 54.180 ;
        RECT 73.310 52.420 73.540 52.430 ;
        RECT 74.560 52.260 75.420 52.650 ;
        RECT 70.400 52.030 75.420 52.260 ;
        RECT 85.140 52.420 85.740 53.030 ;
        RECT 66.660 51.480 69.875 51.710 ;
        RECT 66.660 51.475 67.620 51.480 ;
        RECT 68.540 51.475 69.875 51.480 ;
        RECT 70.420 51.475 71.380 51.705 ;
        RECT 72.300 51.670 73.260 51.705 ;
        RECT 72.300 51.475 73.510 51.670 ;
        RECT 66.280 51.260 66.610 51.270 ;
        RECT 65.790 47.505 66.020 51.025 ;
        RECT 66.280 50.660 66.890 51.260 ;
        RECT 66.380 47.505 66.610 50.660 ;
        RECT 65.790 47.270 66.105 47.505 ;
        RECT 62.900 46.835 63.860 47.065 ;
        RECT 62.960 46.525 63.800 46.835 ;
        RECT 64.065 46.780 64.605 47.270 ;
        RECT 64.055 46.590 64.605 46.780 ;
        RECT 62.900 46.295 63.860 46.525 ;
        RECT 62.535 45.850 62.850 46.090 ;
        RECT 48.770 42.090 49.000 45.850 ;
        RECT 50.025 42.320 50.215 45.850 ;
        RECT 50.650 45.845 50.965 45.850 ;
        RECT 50.650 42.320 50.880 45.845 ;
        RECT 50.020 41.885 50.880 42.320 ;
        RECT 45.880 41.660 46.970 41.870 ;
        RECT 45.880 41.560 46.840 41.660 ;
        RECT 47.760 41.655 48.720 41.885 ;
        RECT 49.640 41.660 50.880 41.885 ;
        RECT 49.640 41.655 50.600 41.660 ;
        RECT 51.380 41.090 52.570 43.250 ;
        RECT 53.040 41.090 54.230 43.250 ;
        RECT 62.620 42.090 62.850 45.850 ;
        RECT 63.285 41.885 63.475 46.295 ;
        RECT 64.065 46.090 64.605 46.590 ;
        RECT 65.915 46.090 66.105 47.270 ;
        RECT 63.910 45.855 64.730 46.090 ;
        RECT 63.910 45.850 64.255 45.855 ;
        RECT 63.910 42.330 64.140 45.850 ;
        RECT 64.500 42.330 64.730 45.855 ;
        RECT 63.910 42.140 64.730 42.330 ;
        RECT 63.910 42.090 64.140 42.140 ;
        RECT 64.500 42.090 64.730 42.140 ;
        RECT 65.790 45.845 66.105 46.090 ;
        RECT 66.275 47.270 66.610 47.505 ;
        RECT 66.275 46.090 66.465 47.270 ;
        RECT 67.045 47.070 67.235 51.475 ;
        RECT 68.920 51.040 69.875 51.475 ;
        RECT 68.925 47.510 69.115 51.040 ;
        RECT 69.550 51.030 69.875 51.040 ;
        RECT 69.550 47.510 69.780 51.030 ;
        RECT 68.925 47.505 69.860 47.510 ;
        RECT 68.925 47.500 69.865 47.505 ;
        RECT 68.920 47.070 69.865 47.500 ;
        RECT 70.805 47.070 70.995 51.475 ;
        RECT 72.680 51.330 73.510 51.475 ;
        RECT 71.240 50.730 71.850 51.330 ;
        RECT 72.680 51.040 73.730 51.330 ;
        RECT 71.430 47.475 71.660 50.730 ;
        RECT 72.685 47.510 72.875 51.040 ;
        RECT 73.120 50.730 73.730 51.040 ;
        RECT 73.310 47.515 73.540 50.730 ;
        RECT 74.100 49.365 74.350 52.030 ;
        RECT 74.870 49.340 76.060 51.500 ;
        RECT 85.140 51.270 85.335 52.420 ;
        RECT 85.945 52.260 86.135 54.580 ;
        RECT 87.440 54.570 88.775 55.350 ;
        RECT 87.825 54.180 88.775 54.570 ;
        RECT 88.955 55.510 89.270 55.765 ;
        RECT 88.955 54.420 89.145 55.510 ;
        RECT 89.705 55.350 89.895 57.670 ;
        RECT 90.330 57.460 90.560 57.510 ;
        RECT 90.920 57.460 91.150 57.510 ;
        RECT 90.330 57.270 91.150 57.460 ;
        RECT 90.330 55.750 90.560 57.270 ;
        RECT 90.920 55.750 91.150 57.270 ;
        RECT 90.330 55.510 91.150 55.750 ;
        RECT 92.210 55.750 92.440 57.510 ;
        RECT 92.210 55.510 92.525 55.750 ;
        RECT 89.320 54.580 90.280 55.350 ;
        RECT 88.955 54.180 89.270 54.420 ;
        RECT 87.825 52.670 88.015 54.180 ;
        RECT 88.450 52.670 88.680 54.180 ;
        RECT 89.040 53.030 89.270 54.180 ;
        RECT 87.820 52.665 88.760 52.670 ;
        RECT 87.820 52.260 88.765 52.665 ;
        RECT 85.560 52.240 86.520 52.260 ;
        RECT 87.440 52.240 88.765 52.260 ;
        RECT 85.560 52.050 88.765 52.240 ;
        RECT 85.560 52.030 86.520 52.050 ;
        RECT 87.440 52.030 88.765 52.050 ;
        RECT 85.560 51.475 86.520 51.705 ;
        RECT 85.140 50.670 85.740 51.270 ;
        RECT 85.280 47.515 85.510 50.670 ;
        RECT 73.310 47.510 73.625 47.515 ;
        RECT 71.430 47.270 71.745 47.475 ;
        RECT 66.660 46.290 67.620 47.070 ;
        RECT 68.540 46.290 69.865 47.070 ;
        RECT 70.400 46.290 71.400 47.070 ;
        RECT 66.275 45.850 66.610 46.090 ;
        RECT 65.790 42.090 66.020 45.845 ;
        RECT 66.380 42.090 66.610 45.850 ;
        RECT 67.045 41.890 67.235 46.290 ;
        RECT 68.925 45.845 69.865 46.290 ;
        RECT 68.925 45.840 69.860 45.845 ;
        RECT 68.925 42.320 69.115 45.840 ;
        RECT 69.550 42.320 69.780 45.840 ;
        RECT 68.925 42.090 69.780 42.320 ;
        RECT 68.925 41.890 69.750 42.090 ;
        RECT 62.900 41.655 63.860 41.885 ;
        RECT 66.660 41.560 67.620 41.890 ;
        RECT 68.540 41.870 69.750 41.890 ;
        RECT 70.805 41.885 70.995 46.290 ;
        RECT 71.555 46.090 71.745 47.270 ;
        RECT 72.685 47.070 73.625 47.510 ;
        RECT 72.280 46.290 73.625 47.070 ;
        RECT 71.430 45.850 71.745 46.090 ;
        RECT 72.685 45.850 73.625 46.290 ;
        RECT 85.195 47.270 85.510 47.515 ;
        RECT 85.195 46.090 85.385 47.270 ;
        RECT 85.945 47.065 86.135 51.475 ;
        RECT 88.575 51.270 88.765 52.030 ;
        RECT 86.570 51.220 86.800 51.270 ;
        RECT 87.160 51.220 87.390 51.270 ;
        RECT 86.570 51.030 87.390 51.220 ;
        RECT 86.570 47.515 86.800 51.030 ;
        RECT 86.570 47.510 86.915 47.515 ;
        RECT 87.160 47.510 87.390 51.030 ;
        RECT 86.570 47.270 87.390 47.510 ;
        RECT 88.450 51.025 88.765 51.270 ;
        RECT 88.940 52.430 89.550 53.030 ;
        RECT 88.940 52.420 89.270 52.430 ;
        RECT 88.940 51.270 89.130 52.420 ;
        RECT 89.705 52.260 89.895 54.580 ;
        RECT 90.465 54.420 91.025 55.510 ;
        RECT 92.335 54.420 92.525 55.510 ;
        RECT 93.465 55.350 93.655 57.670 ;
        RECT 94.090 55.755 94.320 57.510 ;
        RECT 94.090 55.510 94.405 55.755 ;
        RECT 93.060 54.580 94.060 55.350 ;
        RECT 90.330 54.180 91.150 54.420 ;
        RECT 90.330 52.660 90.560 54.180 ;
        RECT 90.920 52.660 91.150 54.180 ;
        RECT 90.330 52.470 91.150 52.660 ;
        RECT 90.330 52.420 90.560 52.470 ;
        RECT 90.920 52.420 91.150 52.470 ;
        RECT 92.210 54.175 92.525 54.420 ;
        RECT 92.210 52.665 92.440 54.175 ;
        RECT 92.210 52.420 92.535 52.665 ;
        RECT 89.320 52.030 90.280 52.260 ;
        RECT 92.345 51.710 92.535 52.420 ;
        RECT 93.465 52.260 93.655 54.580 ;
        RECT 94.215 54.420 94.405 55.510 ;
        RECT 95.345 55.350 95.535 57.670 ;
        RECT 95.970 55.765 96.200 57.510 ;
        RECT 97.220 57.270 98.080 57.670 ;
        RECT 108.250 57.630 109.150 57.670 ;
        RECT 110.130 57.630 111.320 57.670 ;
        RECT 95.970 55.510 96.285 55.765 ;
        RECT 94.940 54.580 95.940 55.350 ;
        RECT 94.090 54.175 94.405 54.420 ;
        RECT 94.090 53.030 94.320 54.175 ;
        RECT 93.910 52.430 94.510 53.030 ;
        RECT 94.090 52.420 94.320 52.430 ;
        RECT 95.345 52.260 95.535 54.580 ;
        RECT 96.095 54.420 96.285 55.510 ;
        RECT 97.220 55.740 97.415 57.270 ;
        RECT 97.850 55.750 98.080 57.270 ;
        RECT 97.850 55.740 98.175 55.750 ;
        RECT 107.940 55.745 108.170 57.510 ;
        RECT 97.220 55.350 98.175 55.740 ;
        RECT 96.820 54.580 98.175 55.350 ;
        RECT 95.970 54.180 96.285 54.420 ;
        RECT 95.970 53.030 96.200 54.180 ;
        RECT 97.220 54.175 98.175 54.580 ;
        RECT 107.855 55.510 108.170 55.745 ;
        RECT 107.855 54.420 108.045 55.510 ;
        RECT 108.605 55.350 108.795 57.630 ;
        RECT 110.480 57.510 111.320 57.630 ;
        RECT 110.480 57.280 111.340 57.510 ;
        RECT 110.485 55.750 110.675 57.280 ;
        RECT 111.110 55.755 111.340 57.280 ;
        RECT 111.700 55.765 111.930 57.510 ;
        RECT 111.110 55.750 111.435 55.755 ;
        RECT 110.485 55.350 111.435 55.750 ;
        RECT 108.220 54.580 109.180 55.350 ;
        RECT 107.855 54.180 108.170 54.420 ;
        RECT 97.220 54.170 98.170 54.175 ;
        RECT 95.790 52.430 96.390 53.030 ;
        RECT 97.220 52.650 97.415 54.170 ;
        RECT 97.850 52.650 98.080 54.170 ;
        RECT 107.940 53.030 108.170 54.180 ;
        RECT 95.970 52.420 96.200 52.430 ;
        RECT 97.220 52.260 98.080 52.650 ;
        RECT 93.060 52.030 98.080 52.260 ;
        RECT 107.800 52.420 108.400 53.030 ;
        RECT 89.320 51.480 92.535 51.710 ;
        RECT 89.320 51.475 90.280 51.480 ;
        RECT 91.200 51.475 92.535 51.480 ;
        RECT 93.080 51.475 94.040 51.705 ;
        RECT 94.960 51.670 95.920 51.705 ;
        RECT 94.960 51.475 96.170 51.670 ;
        RECT 88.940 51.260 89.270 51.270 ;
        RECT 88.450 47.505 88.680 51.025 ;
        RECT 88.940 50.660 89.550 51.260 ;
        RECT 89.040 47.505 89.270 50.660 ;
        RECT 88.450 47.270 88.765 47.505 ;
        RECT 85.560 46.835 86.520 47.065 ;
        RECT 85.620 46.525 86.460 46.835 ;
        RECT 86.725 46.780 87.265 47.270 ;
        RECT 86.715 46.590 87.265 46.780 ;
        RECT 85.560 46.295 86.520 46.525 ;
        RECT 85.195 45.850 85.510 46.090 ;
        RECT 71.430 42.090 71.660 45.850 ;
        RECT 72.685 42.320 72.875 45.850 ;
        RECT 73.310 45.845 73.625 45.850 ;
        RECT 73.310 42.320 73.540 45.845 ;
        RECT 72.680 41.885 73.540 42.320 ;
        RECT 68.540 41.660 69.630 41.870 ;
        RECT 68.540 41.560 69.500 41.660 ;
        RECT 70.420 41.655 71.380 41.885 ;
        RECT 72.300 41.660 73.540 41.885 ;
        RECT 72.300 41.655 73.260 41.660 ;
        RECT 74.040 41.090 75.230 43.250 ;
        RECT 75.700 41.090 76.890 43.250 ;
        RECT 85.280 42.090 85.510 45.850 ;
        RECT 85.945 41.885 86.135 46.295 ;
        RECT 86.725 46.090 87.265 46.590 ;
        RECT 88.575 46.090 88.765 47.270 ;
        RECT 86.570 45.855 87.390 46.090 ;
        RECT 86.570 45.850 86.915 45.855 ;
        RECT 86.570 42.330 86.800 45.850 ;
        RECT 87.160 42.330 87.390 45.855 ;
        RECT 86.570 42.140 87.390 42.330 ;
        RECT 86.570 42.090 86.800 42.140 ;
        RECT 87.160 42.090 87.390 42.140 ;
        RECT 88.450 45.845 88.765 46.090 ;
        RECT 88.935 47.270 89.270 47.505 ;
        RECT 88.935 46.090 89.125 47.270 ;
        RECT 89.705 47.070 89.895 51.475 ;
        RECT 91.580 51.040 92.535 51.475 ;
        RECT 91.585 47.510 91.775 51.040 ;
        RECT 92.210 51.030 92.535 51.040 ;
        RECT 92.210 47.510 92.440 51.030 ;
        RECT 91.585 47.505 92.520 47.510 ;
        RECT 91.585 47.500 92.525 47.505 ;
        RECT 91.580 47.070 92.525 47.500 ;
        RECT 93.465 47.070 93.655 51.475 ;
        RECT 95.340 51.330 96.170 51.475 ;
        RECT 93.900 50.730 94.510 51.330 ;
        RECT 95.340 51.040 96.390 51.330 ;
        RECT 94.090 47.475 94.320 50.730 ;
        RECT 95.345 47.510 95.535 51.040 ;
        RECT 95.780 50.730 96.390 51.040 ;
        RECT 95.970 47.515 96.200 50.730 ;
        RECT 96.760 49.365 97.010 52.030 ;
        RECT 97.530 49.340 98.720 51.500 ;
        RECT 107.800 51.270 107.995 52.420 ;
        RECT 108.605 52.260 108.795 54.580 ;
        RECT 110.100 54.570 111.435 55.350 ;
        RECT 110.485 54.180 111.435 54.570 ;
        RECT 111.615 55.510 111.930 55.765 ;
        RECT 111.615 54.420 111.805 55.510 ;
        RECT 112.365 55.350 112.555 57.670 ;
        RECT 112.990 57.460 113.220 57.510 ;
        RECT 113.580 57.460 113.810 57.510 ;
        RECT 112.990 57.270 113.810 57.460 ;
        RECT 112.990 55.750 113.220 57.270 ;
        RECT 113.580 55.750 113.810 57.270 ;
        RECT 112.990 55.510 113.810 55.750 ;
        RECT 114.870 55.750 115.100 57.510 ;
        RECT 114.870 55.510 115.185 55.750 ;
        RECT 111.980 54.580 112.940 55.350 ;
        RECT 111.615 54.180 111.930 54.420 ;
        RECT 110.485 52.670 110.675 54.180 ;
        RECT 111.110 52.670 111.340 54.180 ;
        RECT 111.700 53.030 111.930 54.180 ;
        RECT 110.480 52.665 111.420 52.670 ;
        RECT 110.480 52.260 111.425 52.665 ;
        RECT 108.220 52.240 109.180 52.260 ;
        RECT 110.100 52.240 111.425 52.260 ;
        RECT 108.220 52.050 111.425 52.240 ;
        RECT 108.220 52.030 109.180 52.050 ;
        RECT 110.100 52.030 111.425 52.050 ;
        RECT 108.220 51.475 109.180 51.705 ;
        RECT 107.800 50.670 108.400 51.270 ;
        RECT 107.940 47.515 108.170 50.670 ;
        RECT 95.970 47.510 96.285 47.515 ;
        RECT 94.090 47.270 94.405 47.475 ;
        RECT 89.320 46.290 90.280 47.070 ;
        RECT 91.200 46.290 92.525 47.070 ;
        RECT 93.060 46.290 94.060 47.070 ;
        RECT 88.935 45.850 89.270 46.090 ;
        RECT 88.450 42.090 88.680 45.845 ;
        RECT 89.040 42.090 89.270 45.850 ;
        RECT 89.705 41.890 89.895 46.290 ;
        RECT 91.585 45.845 92.525 46.290 ;
        RECT 91.585 45.840 92.520 45.845 ;
        RECT 91.585 42.320 91.775 45.840 ;
        RECT 92.210 42.320 92.440 45.840 ;
        RECT 91.585 42.090 92.440 42.320 ;
        RECT 91.585 41.890 92.410 42.090 ;
        RECT 85.560 41.655 86.520 41.885 ;
        RECT 89.320 41.560 90.280 41.890 ;
        RECT 91.200 41.870 92.410 41.890 ;
        RECT 93.465 41.885 93.655 46.290 ;
        RECT 94.215 46.090 94.405 47.270 ;
        RECT 95.345 47.070 96.285 47.510 ;
        RECT 94.940 46.290 96.285 47.070 ;
        RECT 94.090 45.850 94.405 46.090 ;
        RECT 95.345 45.850 96.285 46.290 ;
        RECT 107.855 47.270 108.170 47.515 ;
        RECT 107.855 46.090 108.045 47.270 ;
        RECT 108.605 47.065 108.795 51.475 ;
        RECT 111.235 51.270 111.425 52.030 ;
        RECT 109.230 51.220 109.460 51.270 ;
        RECT 109.820 51.220 110.050 51.270 ;
        RECT 109.230 51.030 110.050 51.220 ;
        RECT 109.230 47.515 109.460 51.030 ;
        RECT 109.230 47.510 109.575 47.515 ;
        RECT 109.820 47.510 110.050 51.030 ;
        RECT 109.230 47.270 110.050 47.510 ;
        RECT 111.110 51.025 111.425 51.270 ;
        RECT 111.600 52.430 112.210 53.030 ;
        RECT 111.600 52.420 111.930 52.430 ;
        RECT 111.600 51.270 111.790 52.420 ;
        RECT 112.365 52.260 112.555 54.580 ;
        RECT 113.125 54.420 113.685 55.510 ;
        RECT 114.995 54.420 115.185 55.510 ;
        RECT 116.125 55.350 116.315 57.670 ;
        RECT 116.750 55.755 116.980 57.510 ;
        RECT 116.750 55.510 117.065 55.755 ;
        RECT 115.720 54.580 116.720 55.350 ;
        RECT 112.990 54.180 113.810 54.420 ;
        RECT 112.990 52.660 113.220 54.180 ;
        RECT 113.580 52.660 113.810 54.180 ;
        RECT 112.990 52.470 113.810 52.660 ;
        RECT 112.990 52.420 113.220 52.470 ;
        RECT 113.580 52.420 113.810 52.470 ;
        RECT 114.870 54.175 115.185 54.420 ;
        RECT 114.870 52.665 115.100 54.175 ;
        RECT 114.870 52.420 115.195 52.665 ;
        RECT 111.980 52.030 112.940 52.260 ;
        RECT 115.005 51.710 115.195 52.420 ;
        RECT 116.125 52.260 116.315 54.580 ;
        RECT 116.875 54.420 117.065 55.510 ;
        RECT 118.005 55.350 118.195 57.670 ;
        RECT 118.630 55.765 118.860 57.510 ;
        RECT 119.880 57.270 120.740 57.670 ;
        RECT 118.630 55.510 118.945 55.765 ;
        RECT 117.600 54.580 118.600 55.350 ;
        RECT 116.750 54.175 117.065 54.420 ;
        RECT 116.750 53.030 116.980 54.175 ;
        RECT 116.570 52.430 117.170 53.030 ;
        RECT 116.750 52.420 116.980 52.430 ;
        RECT 118.005 52.260 118.195 54.580 ;
        RECT 118.755 54.420 118.945 55.510 ;
        RECT 119.880 55.740 120.075 57.270 ;
        RECT 120.510 55.750 120.740 57.270 ;
        RECT 120.510 55.740 120.835 55.750 ;
        RECT 119.880 55.350 120.835 55.740 ;
        RECT 119.480 54.580 120.835 55.350 ;
        RECT 118.630 54.180 118.945 54.420 ;
        RECT 118.630 53.030 118.860 54.180 ;
        RECT 119.880 54.175 120.835 54.580 ;
        RECT 119.880 54.170 120.830 54.175 ;
        RECT 118.450 52.430 119.050 53.030 ;
        RECT 119.880 52.650 120.075 54.170 ;
        RECT 120.510 52.650 120.740 54.170 ;
        RECT 118.630 52.420 118.860 52.430 ;
        RECT 119.880 52.260 120.740 52.650 ;
        RECT 115.720 52.030 120.740 52.260 ;
        RECT 111.980 51.480 115.195 51.710 ;
        RECT 111.980 51.475 112.940 51.480 ;
        RECT 113.860 51.475 115.195 51.480 ;
        RECT 115.740 51.475 116.700 51.705 ;
        RECT 117.620 51.670 118.580 51.705 ;
        RECT 117.620 51.475 118.830 51.670 ;
        RECT 111.600 51.260 111.930 51.270 ;
        RECT 111.110 47.505 111.340 51.025 ;
        RECT 111.600 50.660 112.210 51.260 ;
        RECT 111.700 47.505 111.930 50.660 ;
        RECT 111.110 47.270 111.425 47.505 ;
        RECT 108.220 46.835 109.180 47.065 ;
        RECT 108.280 46.525 109.120 46.835 ;
        RECT 109.385 46.780 109.925 47.270 ;
        RECT 109.375 46.590 109.925 46.780 ;
        RECT 108.220 46.295 109.180 46.525 ;
        RECT 107.855 45.850 108.170 46.090 ;
        RECT 94.090 42.090 94.320 45.850 ;
        RECT 95.345 42.320 95.535 45.850 ;
        RECT 95.970 45.845 96.285 45.850 ;
        RECT 95.970 42.320 96.200 45.845 ;
        RECT 95.340 41.885 96.200 42.320 ;
        RECT 91.200 41.660 92.290 41.870 ;
        RECT 91.200 41.560 92.160 41.660 ;
        RECT 93.080 41.655 94.040 41.885 ;
        RECT 94.960 41.660 96.200 41.885 ;
        RECT 94.960 41.655 95.920 41.660 ;
        RECT 96.700 41.090 97.890 43.250 ;
        RECT 98.360 41.090 99.550 43.250 ;
        RECT 107.940 42.090 108.170 45.850 ;
        RECT 108.605 41.885 108.795 46.295 ;
        RECT 109.385 46.090 109.925 46.590 ;
        RECT 111.235 46.090 111.425 47.270 ;
        RECT 109.230 45.855 110.050 46.090 ;
        RECT 109.230 45.850 109.575 45.855 ;
        RECT 109.230 42.330 109.460 45.850 ;
        RECT 109.820 42.330 110.050 45.855 ;
        RECT 109.230 42.140 110.050 42.330 ;
        RECT 109.230 42.090 109.460 42.140 ;
        RECT 109.820 42.090 110.050 42.140 ;
        RECT 111.110 45.845 111.425 46.090 ;
        RECT 111.595 47.270 111.930 47.505 ;
        RECT 111.595 46.090 111.785 47.270 ;
        RECT 112.365 47.070 112.555 51.475 ;
        RECT 114.240 51.040 115.195 51.475 ;
        RECT 114.245 47.510 114.435 51.040 ;
        RECT 114.870 51.030 115.195 51.040 ;
        RECT 114.870 47.510 115.100 51.030 ;
        RECT 114.245 47.505 115.180 47.510 ;
        RECT 114.245 47.500 115.185 47.505 ;
        RECT 114.240 47.070 115.185 47.500 ;
        RECT 116.125 47.070 116.315 51.475 ;
        RECT 118.000 51.330 118.830 51.475 ;
        RECT 116.560 50.730 117.170 51.330 ;
        RECT 118.000 51.040 119.050 51.330 ;
        RECT 116.750 47.475 116.980 50.730 ;
        RECT 118.005 47.510 118.195 51.040 ;
        RECT 118.440 50.730 119.050 51.040 ;
        RECT 118.630 47.515 118.860 50.730 ;
        RECT 119.420 49.365 119.670 52.030 ;
        RECT 120.190 49.340 121.380 51.500 ;
        RECT 118.630 47.510 118.945 47.515 ;
        RECT 116.750 47.270 117.065 47.475 ;
        RECT 111.980 46.290 112.940 47.070 ;
        RECT 113.860 46.290 115.185 47.070 ;
        RECT 115.720 46.290 116.720 47.070 ;
        RECT 111.595 45.850 111.930 46.090 ;
        RECT 111.110 42.090 111.340 45.845 ;
        RECT 111.700 42.090 111.930 45.850 ;
        RECT 112.365 41.890 112.555 46.290 ;
        RECT 114.245 45.845 115.185 46.290 ;
        RECT 114.245 45.840 115.180 45.845 ;
        RECT 114.245 42.320 114.435 45.840 ;
        RECT 114.870 42.320 115.100 45.840 ;
        RECT 114.245 42.090 115.100 42.320 ;
        RECT 114.245 41.890 115.070 42.090 ;
        RECT 108.220 41.655 109.180 41.885 ;
        RECT 111.980 41.560 112.940 41.890 ;
        RECT 113.860 41.870 115.070 41.890 ;
        RECT 116.125 41.885 116.315 46.290 ;
        RECT 116.875 46.090 117.065 47.270 ;
        RECT 118.005 47.070 118.945 47.510 ;
        RECT 117.600 46.290 118.945 47.070 ;
        RECT 116.750 45.850 117.065 46.090 ;
        RECT 118.005 45.850 118.945 46.290 ;
        RECT 116.750 42.090 116.980 45.850 ;
        RECT 118.005 42.320 118.195 45.850 ;
        RECT 118.630 45.845 118.945 45.850 ;
        RECT 118.630 42.320 118.860 45.845 ;
        RECT 118.000 41.885 118.860 42.320 ;
        RECT 113.860 41.660 114.950 41.870 ;
        RECT 113.860 41.560 114.820 41.660 ;
        RECT 115.740 41.655 116.700 41.885 ;
        RECT 117.620 41.660 118.860 41.885 ;
        RECT 117.620 41.655 118.580 41.660 ;
        RECT 119.360 41.090 120.550 43.250 ;
        RECT 121.020 41.090 122.210 43.250 ;
      LAYER via ;
        RECT 76.380 187.650 76.640 187.910 ;
        RECT 93.400 187.650 93.660 187.910 ;
        RECT 74.540 187.310 74.800 187.570 ;
        RECT 117.320 187.310 117.580 187.570 ;
        RECT 83.740 185.610 84.000 185.870 ;
        RECT 110.420 185.610 110.680 185.870 ;
        RECT 102.140 185.270 102.400 185.530 ;
        RECT 106.740 185.270 107.000 185.530 ;
        RECT 112.260 185.270 112.520 185.530 ;
        RECT 57.060 184.930 57.320 185.190 ;
        RECT 58.440 184.930 58.700 185.190 ;
        RECT 62.580 184.930 62.840 185.190 ;
        RECT 65.800 184.930 66.060 185.190 ;
        RECT 63.960 184.590 64.220 184.850 ;
        RECT 69.940 184.930 70.200 185.190 ;
        RECT 73.160 184.930 73.420 185.190 ;
        RECT 75.920 184.930 76.180 185.190 ;
        RECT 83.280 184.930 83.540 185.190 ;
        RECT 73.620 184.590 73.880 184.850 ;
        RECT 98.460 184.930 98.720 185.190 ;
        RECT 93.860 184.590 94.120 184.850 ;
        RECT 100.760 184.590 101.020 184.850 ;
        RECT 109.960 184.590 110.220 184.850 ;
        RECT 88.800 184.250 89.060 184.510 ;
        RECT 89.260 184.250 89.520 184.510 ;
        RECT 91.100 184.250 91.360 184.510 ;
        RECT 103.060 184.250 103.320 184.510 ;
        RECT 103.980 184.250 104.240 184.510 ;
        RECT 108.120 184.250 108.380 184.510 ;
        RECT 109.500 184.250 109.760 184.510 ;
        RECT 113.180 184.250 113.440 184.510 ;
        RECT 67.180 183.230 67.440 183.490 ;
        RECT 73.160 183.230 73.420 183.490 ;
        RECT 74.540 183.230 74.800 183.490 ;
        RECT 75.000 183.230 75.260 183.490 ;
        RECT 83.740 183.230 84.000 183.490 ;
        RECT 89.260 183.230 89.520 183.490 ;
        RECT 93.860 183.230 94.120 183.490 ;
        RECT 98.460 183.230 98.720 183.490 ;
        RECT 100.300 183.230 100.560 183.490 ;
        RECT 113.180 183.230 113.440 183.490 ;
        RECT 55.220 182.890 55.480 183.150 ;
        RECT 56.600 182.550 56.860 182.810 ;
        RECT 62.120 182.550 62.380 182.810 ;
        RECT 63.500 182.210 63.760 182.470 ;
        RECT 77.300 182.550 77.560 182.810 ;
        RECT 90.640 182.890 90.900 183.150 ;
        RECT 93.400 182.890 93.660 183.150 ;
        RECT 108.120 182.890 108.380 183.150 ;
        RECT 81.900 182.550 82.160 182.810 ;
        RECT 83.280 182.550 83.540 182.810 ;
        RECT 85.580 182.550 85.840 182.810 ;
        RECT 54.300 181.870 54.560 182.130 ;
        RECT 53.840 181.530 54.100 181.790 ;
        RECT 72.700 182.210 72.960 182.470 ;
        RECT 76.380 182.210 76.640 182.470 ;
        RECT 72.700 181.530 72.960 181.790 ;
        RECT 76.840 181.530 77.100 181.790 ;
        RECT 86.040 182.210 86.300 182.470 ;
        RECT 86.500 182.210 86.760 182.470 ;
        RECT 90.180 182.210 90.440 182.470 ;
        RECT 95.700 182.550 95.960 182.810 ;
        RECT 102.600 182.550 102.860 182.810 ;
        RECT 106.740 182.550 107.000 182.810 ;
        RECT 108.580 182.550 108.840 182.810 ;
        RECT 94.780 182.210 95.040 182.470 ;
        RECT 89.720 181.870 89.980 182.130 ;
        RECT 98.920 182.210 99.180 182.470 ;
        RECT 101.680 182.210 101.940 182.470 ;
        RECT 109.040 182.210 109.300 182.470 ;
        RECT 102.140 181.870 102.400 182.130 ;
        RECT 103.520 181.870 103.780 182.130 ;
        RECT 95.240 181.530 95.500 181.790 ;
        RECT 100.300 181.530 100.560 181.790 ;
        RECT 107.660 181.530 107.920 181.790 ;
        RECT 62.580 180.510 62.840 180.770 ;
        RECT 64.880 180.510 65.140 180.770 ;
        RECT 85.580 180.510 85.840 180.770 ;
        RECT 92.020 180.510 92.280 180.770 ;
        RECT 94.780 180.510 95.040 180.770 ;
        RECT 100.760 180.510 101.020 180.770 ;
        RECT 101.680 180.510 101.940 180.770 ;
        RECT 83.280 180.170 83.540 180.430 ;
        RECT 66.260 179.830 66.520 180.090 ;
        RECT 67.180 179.830 67.440 180.090 ;
        RECT 49.700 178.810 49.960 179.070 ;
        RECT 54.300 179.490 54.560 179.750 ;
        RECT 57.520 179.490 57.780 179.750 ;
        RECT 62.580 179.490 62.840 179.750 ;
        RECT 64.880 179.490 65.140 179.750 ;
        RECT 83.740 179.830 84.000 180.090 ;
        RECT 86.500 179.830 86.760 180.090 ;
        RECT 76.840 179.490 77.100 179.750 ;
        RECT 81.900 179.490 82.160 179.750 ;
        RECT 84.660 179.490 84.920 179.750 ;
        RECT 86.040 179.490 86.300 179.750 ;
        RECT 52.460 179.150 52.720 179.410 ;
        RECT 60.280 179.150 60.540 179.410 ;
        RECT 61.200 179.150 61.460 179.410 ;
        RECT 75.460 179.150 75.720 179.410 ;
        RECT 80.060 179.150 80.320 179.410 ;
        RECT 89.720 179.150 89.980 179.410 ;
        RECT 90.180 179.150 90.440 179.410 ;
        RECT 53.840 178.810 54.100 179.070 ;
        RECT 65.340 178.810 65.600 179.070 ;
        RECT 66.720 178.810 66.980 179.070 ;
        RECT 90.640 178.810 90.900 179.070 ;
        RECT 91.560 178.810 91.820 179.070 ;
        RECT 102.140 179.830 102.400 180.090 ;
        RECT 109.500 179.830 109.760 180.090 ;
        RECT 113.640 179.830 113.900 180.090 ;
        RECT 96.160 179.490 96.420 179.750 ;
        RECT 99.840 179.490 100.100 179.750 ;
        RECT 107.660 179.490 107.920 179.750 ;
        RECT 108.580 179.490 108.840 179.750 ;
        RECT 94.320 178.810 94.580 179.070 ;
        RECT 100.300 178.810 100.560 179.070 ;
        RECT 100.760 178.810 101.020 179.070 ;
        RECT 102.600 178.810 102.860 179.070 ;
        RECT 104.440 178.810 104.700 179.070 ;
        RECT 108.580 178.810 108.840 179.070 ;
        RECT 49.700 177.790 49.960 178.050 ;
        RECT 58.440 177.790 58.700 178.050 ;
        RECT 62.120 177.790 62.380 178.050 ;
        RECT 63.500 177.790 63.760 178.050 ;
        RECT 75.920 177.790 76.180 178.050 ;
        RECT 84.200 177.790 84.460 178.050 ;
        RECT 89.260 177.790 89.520 178.050 ;
        RECT 65.340 177.450 65.600 177.710 ;
        RECT 51.540 176.770 51.800 177.030 ;
        RECT 57.520 176.770 57.780 177.030 ;
        RECT 60.740 176.770 61.000 177.030 ;
        RECT 61.200 176.770 61.460 177.030 ;
        RECT 66.260 176.770 66.520 177.030 ;
        RECT 73.160 177.110 73.420 177.370 ;
        RECT 56.600 176.430 56.860 176.690 ;
        RECT 63.500 176.090 63.760 176.350 ;
        RECT 74.080 176.090 74.340 176.350 ;
        RECT 80.060 176.770 80.320 177.030 ;
        RECT 84.200 177.110 84.460 177.370 ;
        RECT 84.660 177.110 84.920 177.370 ;
        RECT 82.360 176.770 82.620 177.030 ;
        RECT 88.800 176.770 89.060 177.030 ;
        RECT 92.020 177.450 92.280 177.710 ;
        RECT 95.240 177.790 95.500 178.050 ;
        RECT 96.620 177.790 96.880 178.050 ;
        RECT 109.960 177.790 110.220 178.050 ;
        RECT 96.160 177.450 96.420 177.710 ;
        RECT 95.240 177.110 95.500 177.370 ;
        RECT 99.380 177.450 99.640 177.710 ;
        RECT 102.140 177.110 102.400 177.370 ;
        RECT 103.520 177.110 103.780 177.370 ;
        RECT 104.900 177.110 105.160 177.370 ;
        RECT 112.260 177.110 112.520 177.370 ;
        RECT 96.620 176.770 96.880 177.030 ;
        RECT 99.840 176.770 100.100 177.030 ;
        RECT 100.300 176.770 100.560 177.030 ;
        RECT 104.440 176.770 104.700 177.030 ;
        RECT 92.940 176.430 93.200 176.690 ;
        RECT 89.260 176.090 89.520 176.350 ;
        RECT 93.400 176.090 93.660 176.350 ;
        RECT 99.380 176.090 99.640 176.350 ;
        RECT 103.060 176.090 103.320 176.350 ;
        RECT 104.440 176.090 104.700 176.350 ;
        RECT 111.340 176.770 111.600 177.030 ;
        RECT 60.740 175.070 61.000 175.330 ;
        RECT 52.460 174.390 52.720 174.650 ;
        RECT 61.200 174.390 61.460 174.650 ;
        RECT 72.700 174.730 72.960 174.990 ;
        RECT 74.080 174.730 74.340 174.990 ;
        RECT 86.040 175.070 86.300 175.330 ;
        RECT 89.720 175.070 89.980 175.330 ;
        RECT 93.400 175.070 93.660 175.330 ;
        RECT 96.620 175.070 96.880 175.330 ;
        RECT 84.660 174.730 84.920 174.990 ;
        RECT 52.000 174.050 52.260 174.310 ;
        RECT 55.220 174.050 55.480 174.310 ;
        RECT 58.900 174.050 59.160 174.310 ;
        RECT 59.360 174.050 59.620 174.310 ;
        RECT 67.640 174.050 67.900 174.310 ;
        RECT 82.820 174.390 83.080 174.650 ;
        RECT 69.940 174.050 70.200 174.310 ;
        RECT 72.240 174.050 72.500 174.310 ;
        RECT 75.000 174.050 75.260 174.310 ;
        RECT 76.380 174.050 76.640 174.310 ;
        RECT 84.660 174.050 84.920 174.310 ;
        RECT 89.260 174.390 89.520 174.650 ;
        RECT 99.840 174.390 100.100 174.650 ;
        RECT 90.180 174.050 90.440 174.310 ;
        RECT 94.320 174.050 94.580 174.310 ;
        RECT 101.680 174.390 101.940 174.650 ;
        RECT 102.600 174.390 102.860 174.650 ;
        RECT 103.060 174.390 103.320 174.650 ;
        RECT 104.440 174.390 104.700 174.650 ;
        RECT 56.140 173.370 56.400 173.630 ;
        RECT 58.440 173.370 58.700 173.630 ;
        RECT 63.500 173.370 63.760 173.630 ;
        RECT 65.800 173.370 66.060 173.630 ;
        RECT 66.260 173.370 66.520 173.630 ;
        RECT 68.100 173.370 68.360 173.630 ;
        RECT 75.000 173.370 75.260 173.630 ;
        RECT 76.380 173.370 76.640 173.630 ;
        RECT 85.120 173.370 85.380 173.630 ;
        RECT 86.040 173.370 86.300 173.630 ;
        RECT 87.880 173.370 88.140 173.630 ;
        RECT 93.860 173.370 94.120 173.630 ;
        RECT 94.320 173.370 94.580 173.630 ;
        RECT 98.460 173.710 98.720 173.970 ;
        RECT 109.500 174.390 109.760 174.650 ;
        RECT 112.260 174.390 112.520 174.650 ;
        RECT 108.580 174.050 108.840 174.310 ;
        RECT 109.040 174.050 109.300 174.310 ;
        RECT 105.820 173.710 106.080 173.970 ;
        RECT 99.840 173.370 100.100 173.630 ;
        RECT 100.300 173.370 100.560 173.630 ;
        RECT 104.900 173.370 105.160 173.630 ;
        RECT 111.800 173.370 112.060 173.630 ;
        RECT 113.180 173.370 113.440 173.630 ;
        RECT 114.560 173.370 114.820 173.630 ;
        RECT 57.060 172.350 57.320 172.610 ;
        RECT 44.640 171.670 44.900 171.930 ;
        RECT 68.100 172.350 68.360 172.610 ;
        RECT 72.240 172.350 72.500 172.610 ;
        RECT 83.280 172.350 83.540 172.610 ;
        RECT 88.340 172.350 88.600 172.610 ;
        RECT 89.260 172.350 89.520 172.610 ;
        RECT 94.780 172.350 95.040 172.610 ;
        RECT 98.000 172.350 98.260 172.610 ;
        RECT 103.980 172.350 104.240 172.610 ;
        RECT 64.420 172.010 64.680 172.270 ;
        RECT 58.900 171.670 59.160 171.930 ;
        RECT 54.300 171.330 54.560 171.590 ;
        RECT 60.740 171.330 61.000 171.590 ;
        RECT 65.800 171.670 66.060 171.930 ;
        RECT 66.260 171.670 66.520 171.930 ;
        RECT 69.940 172.010 70.200 172.270 ;
        RECT 72.700 172.010 72.960 172.270 ;
        RECT 75.920 172.010 76.180 172.270 ;
        RECT 87.420 172.010 87.680 172.270 ;
        RECT 82.820 171.670 83.080 171.930 ;
        RECT 86.960 171.670 87.220 171.930 ;
        RECT 101.680 172.010 101.940 172.270 ;
        RECT 104.440 172.010 104.700 172.270 ;
        RECT 98.460 171.670 98.720 171.930 ;
        RECT 98.920 171.670 99.180 171.930 ;
        RECT 104.900 171.670 105.160 171.930 ;
        RECT 108.580 172.350 108.840 172.610 ;
        RECT 109.500 171.670 109.760 171.930 ;
        RECT 66.720 171.330 66.980 171.590 ;
        RECT 87.880 170.990 88.140 171.250 ;
        RECT 95.240 171.330 95.500 171.590 ;
        RECT 94.780 170.990 95.040 171.250 ;
        RECT 99.840 170.990 100.100 171.250 ;
        RECT 100.300 170.990 100.560 171.250 ;
        RECT 54.760 170.650 55.020 170.910 ;
        RECT 68.100 170.650 68.360 170.910 ;
        RECT 80.980 170.650 81.240 170.910 ;
        RECT 81.440 170.650 81.700 170.910 ;
        RECT 87.420 170.650 87.680 170.910 ;
        RECT 93.860 170.650 94.120 170.910 ;
        RECT 104.900 170.650 105.160 170.910 ;
        RECT 105.820 170.650 106.080 170.910 ;
        RECT 109.960 170.650 110.220 170.910 ;
        RECT 63.960 169.630 64.220 169.890 ;
        RECT 75.920 169.630 76.180 169.890 ;
        RECT 83.280 169.630 83.540 169.890 ;
        RECT 74.080 169.290 74.340 169.550 ;
        RECT 60.740 168.950 61.000 169.210 ;
        RECT 67.640 168.950 67.900 169.210 ;
        RECT 55.220 168.610 55.480 168.870 ;
        RECT 68.100 168.610 68.360 168.870 ;
        RECT 68.560 168.610 68.820 168.870 ;
        RECT 72.700 168.950 72.960 169.210 ;
        RECT 81.440 168.950 81.700 169.210 ;
        RECT 83.740 168.950 84.000 169.210 ;
        RECT 90.180 169.630 90.440 169.890 ;
        RECT 98.920 169.630 99.180 169.890 ;
        RECT 103.520 169.630 103.780 169.890 ;
        RECT 57.980 167.930 58.240 168.190 ;
        RECT 64.420 168.270 64.680 168.530 ;
        RECT 76.840 168.270 77.100 168.530 ;
        RECT 81.440 168.270 81.700 168.530 ;
        RECT 71.780 167.930 72.040 168.190 ;
        RECT 82.820 168.610 83.080 168.870 ;
        RECT 86.960 168.950 87.220 169.210 ;
        RECT 94.320 169.290 94.580 169.550 ;
        RECT 104.900 169.290 105.160 169.550 ;
        RECT 95.700 168.950 95.960 169.210 ;
        RECT 98.000 168.950 98.260 169.210 ;
        RECT 100.300 168.950 100.560 169.210 ;
        RECT 101.220 168.950 101.480 169.210 ;
        RECT 112.260 169.290 112.520 169.550 ;
        RECT 109.500 168.950 109.760 169.210 ;
        RECT 87.880 168.610 88.140 168.870 ;
        RECT 93.400 168.610 93.660 168.870 ;
        RECT 93.860 168.610 94.120 168.870 ;
        RECT 90.180 167.930 90.440 168.190 ;
        RECT 92.940 167.930 93.200 168.190 ;
        RECT 101.680 168.610 101.940 168.870 ;
        RECT 102.600 168.610 102.860 168.870 ;
        RECT 100.300 167.930 100.560 168.190 ;
        RECT 102.600 167.930 102.860 168.190 ;
        RECT 108.120 167.930 108.380 168.190 ;
        RECT 109.960 167.930 110.220 168.190 ;
        RECT 54.300 166.910 54.560 167.170 ;
        RECT 54.760 166.910 55.020 167.170 ;
        RECT 54.760 166.230 55.020 166.490 ;
        RECT 55.220 166.230 55.480 166.490 ;
        RECT 68.560 166.910 68.820 167.170 ;
        RECT 71.780 166.570 72.040 166.830 ;
        RECT 77.760 166.570 78.020 166.830 ;
        RECT 75.460 166.230 75.720 166.490 ;
        RECT 93.400 166.910 93.660 167.170 ;
        RECT 102.600 166.910 102.860 167.170 ;
        RECT 103.980 166.910 104.240 167.170 ;
        RECT 109.500 166.910 109.760 167.170 ;
        RECT 80.520 166.570 80.780 166.830 ;
        RECT 81.440 166.230 81.700 166.490 ;
        RECT 92.020 166.230 92.280 166.490 ;
        RECT 92.480 166.230 92.740 166.490 ;
        RECT 93.860 166.230 94.120 166.490 ;
        RECT 111.800 166.570 112.060 166.830 ;
        RECT 53.840 165.890 54.100 166.150 ;
        RECT 58.440 165.890 58.700 166.150 ;
        RECT 59.820 165.890 60.080 166.150 ;
        RECT 57.520 165.550 57.780 165.810 ;
        RECT 59.820 165.210 60.080 165.470 ;
        RECT 72.700 165.210 72.960 165.470 ;
        RECT 96.160 166.230 96.420 166.490 ;
        RECT 101.680 166.230 101.940 166.490 ;
        RECT 103.980 166.230 104.240 166.490 ;
        RECT 104.440 165.890 104.700 166.150 ;
        RECT 105.360 166.230 105.620 166.490 ;
        RECT 110.880 166.230 111.140 166.490 ;
        RECT 108.120 165.890 108.380 166.150 ;
        RECT 103.520 165.550 103.780 165.810 ;
        RECT 111.340 165.550 111.600 165.810 ;
        RECT 96.620 165.210 96.880 165.470 ;
        RECT 109.960 165.210 110.220 165.470 ;
        RECT 63.500 164.190 63.760 164.450 ;
        RECT 55.220 163.510 55.480 163.770 ;
        RECT 82.360 164.190 82.620 164.450 ;
        RECT 86.500 164.190 86.760 164.450 ;
        RECT 92.480 164.190 92.740 164.450 ;
        RECT 96.620 164.190 96.880 164.450 ;
        RECT 103.060 164.190 103.320 164.450 ;
        RECT 116.860 164.190 117.120 164.450 ;
        RECT 67.180 163.850 67.440 164.110 ;
        RECT 70.860 163.850 71.120 164.110 ;
        RECT 75.000 163.850 75.260 164.110 ;
        RECT 82.820 163.850 83.080 164.110 ;
        RECT 59.820 163.170 60.080 163.430 ;
        RECT 53.840 162.830 54.100 163.090 ;
        RECT 69.480 163.510 69.740 163.770 ;
        RECT 73.160 163.510 73.420 163.770 ;
        RECT 65.340 163.170 65.600 163.430 ;
        RECT 65.800 163.170 66.060 163.430 ;
        RECT 69.940 163.170 70.200 163.430 ;
        RECT 72.700 163.170 72.960 163.430 ;
        RECT 55.220 162.490 55.480 162.750 ;
        RECT 65.340 162.490 65.600 162.750 ;
        RECT 77.760 162.490 78.020 162.750 ;
        RECT 81.440 163.170 81.700 163.430 ;
        RECT 82.360 163.170 82.620 163.430 ;
        RECT 85.120 163.170 85.380 163.430 ;
        RECT 89.720 163.510 89.980 163.770 ;
        RECT 90.180 163.510 90.440 163.770 ;
        RECT 94.780 163.510 95.040 163.770 ;
        RECT 104.440 163.850 104.700 164.110 ;
        RECT 105.820 163.850 106.080 164.110 ;
        RECT 107.200 163.850 107.460 164.110 ;
        RECT 101.220 163.510 101.480 163.770 ;
        RECT 95.240 163.170 95.500 163.430 ;
        RECT 109.960 163.170 110.220 163.430 ;
        RECT 89.260 162.830 89.520 163.090 ;
        RECT 101.220 162.830 101.480 163.090 ;
        RECT 102.600 162.830 102.860 163.090 ;
        RECT 103.980 162.830 104.240 163.090 ;
        RECT 96.160 162.490 96.420 162.750 ;
        RECT 98.460 162.490 98.720 162.750 ;
        RECT 99.380 162.490 99.640 162.750 ;
        RECT 109.040 162.490 109.300 162.750 ;
        RECT 54.760 161.470 55.020 161.730 ;
        RECT 57.980 161.470 58.240 161.730 ;
        RECT 52.920 160.790 53.180 161.050 ;
        RECT 65.340 161.470 65.600 161.730 ;
        RECT 70.400 161.470 70.660 161.730 ;
        RECT 73.620 161.470 73.880 161.730 ;
        RECT 76.380 161.470 76.640 161.730 ;
        RECT 98.460 161.470 98.720 161.730 ;
        RECT 102.600 161.470 102.860 161.730 ;
        RECT 103.060 161.470 103.320 161.730 ;
        RECT 55.220 160.450 55.480 160.710 ;
        RECT 65.800 161.130 66.060 161.390 ;
        RECT 76.840 161.130 77.100 161.390 ;
        RECT 69.480 160.790 69.740 161.050 ;
        RECT 75.000 160.790 75.260 161.050 ;
        RECT 69.940 160.450 70.200 160.710 ;
        RECT 72.240 160.450 72.500 160.710 ;
        RECT 74.080 160.450 74.340 160.710 ;
        RECT 76.380 160.450 76.640 160.710 ;
        RECT 100.300 161.130 100.560 161.390 ;
        RECT 103.980 161.130 104.240 161.390 ;
        RECT 105.360 161.470 105.620 161.730 ;
        RECT 110.880 161.470 111.140 161.730 ;
        RECT 112.260 161.470 112.520 161.730 ;
        RECT 82.360 160.790 82.620 161.050 ;
        RECT 91.560 160.790 91.820 161.050 ;
        RECT 67.640 160.110 67.900 160.370 ;
        RECT 92.020 160.450 92.280 160.710 ;
        RECT 96.160 160.450 96.420 160.710 ;
        RECT 104.440 160.450 104.700 160.710 ;
        RECT 104.900 160.450 105.160 160.710 ;
        RECT 108.580 160.110 108.840 160.370 ;
        RECT 67.180 159.770 67.440 160.030 ;
        RECT 80.980 159.770 81.240 160.030 ;
        RECT 81.440 159.770 81.700 160.030 ;
        RECT 89.720 159.770 89.980 160.030 ;
        RECT 44.640 158.750 44.900 159.010 ;
        RECT 56.140 158.750 56.400 159.010 ;
        RECT 61.660 158.750 61.920 159.010 ;
        RECT 64.420 158.750 64.680 159.010 ;
        RECT 67.180 158.750 67.440 159.010 ;
        RECT 67.640 158.750 67.900 159.010 ;
        RECT 72.240 158.750 72.500 159.010 ;
        RECT 75.000 158.750 75.260 159.010 ;
        RECT 77.300 158.750 77.560 159.010 ;
        RECT 81.440 158.750 81.700 159.010 ;
        RECT 89.260 158.750 89.520 159.010 ;
        RECT 89.720 158.750 89.980 159.010 ;
        RECT 90.640 158.750 90.900 159.010 ;
        RECT 95.700 158.750 95.960 159.010 ;
        RECT 100.760 158.750 101.020 159.010 ;
        RECT 101.220 158.750 101.480 159.010 ;
        RECT 108.120 158.750 108.380 159.010 ;
        RECT 111.800 158.750 112.060 159.010 ;
        RECT 62.580 158.410 62.840 158.670 ;
        RECT 52.920 158.070 53.180 158.330 ;
        RECT 43.720 157.730 43.980 157.990 ;
        RECT 48.780 157.730 49.040 157.990 ;
        RECT 53.380 157.730 53.640 157.990 ;
        RECT 58.900 157.730 59.160 157.990 ;
        RECT 63.960 157.730 64.220 157.990 ;
        RECT 69.940 157.730 70.200 157.990 ;
        RECT 80.980 158.070 81.240 158.330 ;
        RECT 108.580 158.410 108.840 158.670 ;
        RECT 74.080 157.730 74.340 157.990 ;
        RECT 75.920 157.730 76.180 157.990 ;
        RECT 76.380 157.730 76.640 157.990 ;
        RECT 80.060 157.730 80.320 157.990 ;
        RECT 83.740 157.390 84.000 157.650 ;
        RECT 89.260 157.730 89.520 157.990 ;
        RECT 91.560 157.730 91.820 157.990 ;
        RECT 94.320 157.730 94.580 157.990 ;
        RECT 99.380 157.730 99.640 157.990 ;
        RECT 104.440 157.730 104.700 157.990 ;
        RECT 107.660 157.730 107.920 157.990 ;
        RECT 109.040 157.730 109.300 157.990 ;
        RECT 114.100 157.730 114.360 157.990 ;
        RECT 113.640 157.390 113.900 157.650 ;
        RECT 114.560 157.050 114.820 157.310 ;
        RECT 79.140 156.030 79.400 156.290 ;
        RECT 80.060 156.030 80.320 156.290 ;
        RECT 78.940 128.340 79.200 128.600 ;
        RECT 101.585 128.340 101.845 128.600 ;
        RECT 62.960 127.680 63.800 127.940 ;
        RECT 64.840 127.680 65.680 127.940 ;
        RECT 70.480 127.720 71.320 127.980 ;
        RECT 72.360 127.720 73.200 127.980 ;
        RECT 74.240 127.720 75.080 127.980 ;
        RECT 62.960 124.630 63.800 125.340 ;
        RECT 64.840 124.630 65.680 125.340 ;
        RECT 60.690 123.190 60.960 124.190 ;
        RECT 62.520 122.480 63.030 123.000 ;
        RECT 57.540 120.320 58.460 121.240 ;
        RECT 66.720 124.630 67.560 125.340 ;
        RECT 61.290 120.320 62.210 121.240 ;
        RECT 62.520 120.730 63.030 121.250 ;
        RECT 62.960 116.345 63.800 117.055 ;
        RECT 64.100 115.910 64.570 117.490 ;
        RECT 66.330 122.500 66.840 123.010 ;
        RECT 67.885 124.290 68.285 125.690 ;
        RECT 68.600 124.630 69.440 125.340 ;
        RECT 70.480 124.630 71.320 125.340 ;
        RECT 85.620 127.680 86.460 127.940 ;
        RECT 87.500 127.680 88.340 127.940 ;
        RECT 93.140 127.720 93.980 127.980 ;
        RECT 95.020 127.720 95.860 127.980 ;
        RECT 96.900 127.720 97.740 127.980 ;
        RECT 72.360 124.630 73.200 125.340 ;
        RECT 71.300 122.500 71.800 123.000 ;
        RECT 74.240 124.630 75.080 125.340 ;
        RECT 76.120 124.720 76.670 125.170 ;
        RECT 77.700 124.810 77.960 125.070 ;
        RECT 78.880 124.620 79.230 126.780 ;
        RECT 85.620 124.630 86.460 125.340 ;
        RECT 87.500 124.630 88.340 125.340 ;
        RECT 73.180 122.500 73.680 123.000 ;
        RECT 66.330 120.720 66.840 121.240 ;
        RECT 64.840 116.345 65.680 117.055 ;
        RECT 71.300 120.800 71.800 121.300 ;
        RECT 73.180 120.800 73.680 121.300 ;
        RECT 78.880 120.120 79.230 122.280 ;
        RECT 81.550 123.190 81.820 124.190 ;
        RECT 85.180 122.480 85.690 123.000 ;
        RECT 80.200 120.320 81.120 121.240 ;
        RECT 89.380 124.630 90.220 125.340 ;
        RECT 83.950 120.320 84.870 121.240 ;
        RECT 85.180 120.730 85.690 121.250 ;
        RECT 66.720 116.345 67.560 117.055 ;
        RECT 68.600 116.345 69.440 117.055 ;
        RECT 70.480 116.340 71.320 117.060 ;
        RECT 66.720 111.615 67.560 111.875 ;
        RECT 72.360 116.340 73.200 117.060 ;
        RECT 78.880 116.830 79.230 118.990 ;
        RECT 85.620 116.345 86.460 117.055 ;
        RECT 68.600 111.615 69.440 111.875 ;
        RECT 78.880 112.330 79.230 114.490 ;
        RECT 86.760 115.910 87.230 117.490 ;
        RECT 88.990 122.500 89.500 123.010 ;
        RECT 90.545 124.290 90.945 125.690 ;
        RECT 91.260 124.630 92.100 125.340 ;
        RECT 93.140 124.630 93.980 125.340 ;
        RECT 108.280 127.680 109.120 127.940 ;
        RECT 110.160 127.680 111.000 127.940 ;
        RECT 115.800 127.720 116.640 127.980 ;
        RECT 117.680 127.720 118.520 127.980 ;
        RECT 119.560 127.720 120.400 127.980 ;
        RECT 95.020 124.630 95.860 125.340 ;
        RECT 93.960 122.500 94.460 123.000 ;
        RECT 96.900 124.630 97.740 125.340 ;
        RECT 98.780 124.720 99.330 125.170 ;
        RECT 100.360 124.810 100.620 125.070 ;
        RECT 101.540 124.620 101.890 126.780 ;
        RECT 108.280 124.630 109.120 125.340 ;
        RECT 110.160 124.630 111.000 125.340 ;
        RECT 95.840 122.500 96.340 123.000 ;
        RECT 88.990 120.720 89.500 121.240 ;
        RECT 87.500 116.345 88.340 117.055 ;
        RECT 93.960 120.800 94.460 121.300 ;
        RECT 95.840 120.800 96.340 121.300 ;
        RECT 101.540 120.120 101.890 122.280 ;
        RECT 106.010 123.190 106.280 124.190 ;
        RECT 107.840 122.480 108.350 123.000 ;
        RECT 102.860 120.320 103.780 121.240 ;
        RECT 112.040 124.630 112.880 125.340 ;
        RECT 106.610 120.320 107.530 121.240 ;
        RECT 107.840 120.730 108.350 121.250 ;
        RECT 89.380 116.345 90.220 117.055 ;
        RECT 91.260 116.345 92.100 117.055 ;
        RECT 93.140 116.340 93.980 117.060 ;
        RECT 89.380 111.615 90.220 111.875 ;
        RECT 95.020 116.340 95.860 117.060 ;
        RECT 101.540 116.830 101.890 118.990 ;
        RECT 108.280 116.345 109.120 117.055 ;
        RECT 91.260 111.615 92.100 111.875 ;
        RECT 101.540 112.330 101.890 114.490 ;
        RECT 109.420 115.910 109.890 117.490 ;
        RECT 111.650 122.500 112.160 123.010 ;
        RECT 113.205 124.290 113.605 125.690 ;
        RECT 113.920 124.630 114.760 125.340 ;
        RECT 115.800 124.630 116.640 125.340 ;
        RECT 117.680 124.630 118.520 125.340 ;
        RECT 116.620 122.500 117.120 123.000 ;
        RECT 119.560 124.630 120.400 125.340 ;
        RECT 121.440 124.720 121.990 125.170 ;
        RECT 123.020 124.810 123.280 125.070 ;
        RECT 118.500 122.500 119.000 123.000 ;
        RECT 111.650 120.720 112.160 121.240 ;
        RECT 110.160 116.345 111.000 117.055 ;
        RECT 116.620 120.800 117.120 121.300 ;
        RECT 118.500 120.800 119.000 121.300 ;
        RECT 124.200 120.120 124.550 122.280 ;
        RECT 112.040 116.345 112.880 117.055 ;
        RECT 113.920 116.345 114.760 117.055 ;
        RECT 115.800 116.340 116.640 117.060 ;
        RECT 112.040 111.615 112.880 111.875 ;
        RECT 117.680 116.340 118.520 117.060 ;
        RECT 124.200 116.830 124.550 118.990 ;
        RECT 113.920 111.615 114.760 111.875 ;
        RECT 124.200 112.330 124.550 114.490 ;
        RECT 40.300 110.340 41.140 110.600 ;
        RECT 42.180 110.340 43.020 110.600 ;
        RECT 47.820 110.380 48.660 110.640 ;
        RECT 49.700 110.380 50.540 110.640 ;
        RECT 51.580 110.380 52.420 110.640 ;
        RECT 40.300 107.290 41.140 108.000 ;
        RECT 42.180 107.290 43.020 108.000 ;
        RECT 36.830 105.850 37.100 106.850 ;
        RECT 39.860 105.140 40.370 105.660 ;
        RECT 34.880 102.980 35.800 103.900 ;
        RECT 44.060 107.290 44.900 108.000 ;
        RECT 38.630 102.980 39.550 103.900 ;
        RECT 39.860 103.390 40.370 103.910 ;
        RECT 40.300 99.005 41.140 99.715 ;
        RECT 41.440 98.570 41.910 100.150 ;
        RECT 43.670 105.160 44.180 105.670 ;
        RECT 45.225 106.950 45.625 108.350 ;
        RECT 45.940 107.290 46.780 108.000 ;
        RECT 47.820 107.290 48.660 108.000 ;
        RECT 62.960 110.340 63.800 110.600 ;
        RECT 64.840 110.340 65.680 110.600 ;
        RECT 70.480 110.380 71.320 110.640 ;
        RECT 72.360 110.380 73.200 110.640 ;
        RECT 74.240 110.380 75.080 110.640 ;
        RECT 49.700 107.290 50.540 108.000 ;
        RECT 48.640 105.160 49.140 105.660 ;
        RECT 51.580 107.290 52.420 108.000 ;
        RECT 53.460 107.380 54.010 107.830 ;
        RECT 55.040 107.470 55.300 107.730 ;
        RECT 62.960 107.290 63.800 108.000 ;
        RECT 64.840 107.290 65.680 108.000 ;
        RECT 50.520 105.160 51.020 105.660 ;
        RECT 43.670 103.380 44.180 103.900 ;
        RECT 42.180 99.005 43.020 99.715 ;
        RECT 48.640 103.460 49.140 103.960 ;
        RECT 50.520 103.460 51.020 103.960 ;
        RECT 56.220 102.780 56.570 104.940 ;
        RECT 60.090 105.850 60.360 106.850 ;
        RECT 62.520 105.140 63.030 105.660 ;
        RECT 57.540 102.980 58.460 103.900 ;
        RECT 66.720 107.290 67.560 108.000 ;
        RECT 61.290 102.980 62.210 103.900 ;
        RECT 62.520 103.390 63.030 103.910 ;
        RECT 44.060 99.005 44.900 99.715 ;
        RECT 45.940 99.005 46.780 99.715 ;
        RECT 47.820 99.000 48.660 99.720 ;
        RECT 44.060 94.275 44.900 94.535 ;
        RECT 49.700 99.000 50.540 99.720 ;
        RECT 56.220 99.490 56.570 101.650 ;
        RECT 62.960 99.005 63.800 99.715 ;
        RECT 45.940 94.275 46.780 94.535 ;
        RECT 56.220 94.990 56.570 97.150 ;
        RECT 64.100 98.570 64.570 100.150 ;
        RECT 66.330 105.160 66.840 105.670 ;
        RECT 67.885 106.950 68.285 108.350 ;
        RECT 68.600 107.290 69.440 108.000 ;
        RECT 70.480 107.290 71.320 108.000 ;
        RECT 85.620 110.340 86.460 110.600 ;
        RECT 87.500 110.340 88.340 110.600 ;
        RECT 93.140 110.380 93.980 110.640 ;
        RECT 95.020 110.380 95.860 110.640 ;
        RECT 96.900 110.380 97.740 110.640 ;
        RECT 72.360 107.290 73.200 108.000 ;
        RECT 71.300 105.160 71.800 105.660 ;
        RECT 74.240 107.290 75.080 108.000 ;
        RECT 76.120 107.380 76.670 107.830 ;
        RECT 77.700 107.470 77.960 107.730 ;
        RECT 78.880 107.280 79.230 109.440 ;
        RECT 85.620 107.290 86.460 108.000 ;
        RECT 87.500 107.290 88.340 108.000 ;
        RECT 73.180 105.160 73.680 105.660 ;
        RECT 66.330 103.380 66.840 103.900 ;
        RECT 64.840 99.005 65.680 99.715 ;
        RECT 71.300 103.460 71.800 103.960 ;
        RECT 73.180 103.460 73.680 103.960 ;
        RECT 78.880 102.780 79.230 104.940 ;
        RECT 82.150 105.850 82.420 106.850 ;
        RECT 85.180 105.140 85.690 105.660 ;
        RECT 80.200 102.980 81.120 103.900 ;
        RECT 89.380 107.290 90.220 108.000 ;
        RECT 83.950 102.980 84.870 103.900 ;
        RECT 85.180 103.390 85.690 103.910 ;
        RECT 66.720 99.005 67.560 99.715 ;
        RECT 68.600 99.005 69.440 99.715 ;
        RECT 70.480 99.000 71.320 99.720 ;
        RECT 66.720 94.275 67.560 94.535 ;
        RECT 72.360 99.000 73.200 99.720 ;
        RECT 78.880 99.490 79.230 101.650 ;
        RECT 85.620 99.005 86.460 99.715 ;
        RECT 68.600 94.275 69.440 94.535 ;
        RECT 78.880 94.990 79.230 97.150 ;
        RECT 86.760 98.570 87.230 100.150 ;
        RECT 88.990 105.160 89.500 105.670 ;
        RECT 90.545 106.950 90.945 108.350 ;
        RECT 91.260 107.290 92.100 108.000 ;
        RECT 93.140 107.290 93.980 108.000 ;
        RECT 108.280 110.340 109.120 110.600 ;
        RECT 110.160 110.340 111.000 110.600 ;
        RECT 115.800 110.380 116.640 110.640 ;
        RECT 117.680 110.380 118.520 110.640 ;
        RECT 119.560 110.380 120.400 110.640 ;
        RECT 95.020 107.290 95.860 108.000 ;
        RECT 93.960 105.160 94.460 105.660 ;
        RECT 96.900 107.290 97.740 108.000 ;
        RECT 98.780 107.380 99.330 107.830 ;
        RECT 100.360 107.470 100.620 107.730 ;
        RECT 101.540 107.280 101.890 109.440 ;
        RECT 108.280 107.290 109.120 108.000 ;
        RECT 110.160 107.290 111.000 108.000 ;
        RECT 95.840 105.160 96.340 105.660 ;
        RECT 88.990 103.380 89.500 103.900 ;
        RECT 87.500 99.005 88.340 99.715 ;
        RECT 93.960 103.460 94.460 103.960 ;
        RECT 95.840 103.460 96.340 103.960 ;
        RECT 101.540 102.780 101.890 104.940 ;
        RECT 105.410 105.850 105.680 106.850 ;
        RECT 107.840 105.140 108.350 105.660 ;
        RECT 102.860 102.980 103.780 103.900 ;
        RECT 112.040 107.290 112.880 108.000 ;
        RECT 106.610 102.980 107.530 103.900 ;
        RECT 107.840 103.390 108.350 103.910 ;
        RECT 89.380 99.005 90.220 99.715 ;
        RECT 91.260 99.005 92.100 99.715 ;
        RECT 93.140 99.000 93.980 99.720 ;
        RECT 89.380 94.275 90.220 94.535 ;
        RECT 95.020 99.000 95.860 99.720 ;
        RECT 101.540 99.490 101.890 101.650 ;
        RECT 108.280 99.005 109.120 99.715 ;
        RECT 91.260 94.275 92.100 94.535 ;
        RECT 101.540 94.990 101.890 97.150 ;
        RECT 109.420 98.570 109.890 100.150 ;
        RECT 111.650 105.160 112.160 105.670 ;
        RECT 113.205 106.950 113.605 108.350 ;
        RECT 113.920 107.290 114.760 108.000 ;
        RECT 115.800 107.290 116.640 108.000 ;
        RECT 117.680 107.290 118.520 108.000 ;
        RECT 116.620 105.160 117.120 105.660 ;
        RECT 119.560 107.290 120.400 108.000 ;
        RECT 121.440 107.380 121.990 107.830 ;
        RECT 123.020 107.470 123.280 107.730 ;
        RECT 124.200 107.280 124.550 109.440 ;
        RECT 118.500 105.160 119.000 105.660 ;
        RECT 111.650 103.380 112.160 103.900 ;
        RECT 110.160 99.005 111.000 99.715 ;
        RECT 116.620 103.460 117.120 103.960 ;
        RECT 118.500 103.460 119.000 103.960 ;
        RECT 124.200 102.780 124.550 104.940 ;
        RECT 112.040 99.005 112.880 99.715 ;
        RECT 113.920 99.005 114.760 99.715 ;
        RECT 115.800 99.000 116.640 99.720 ;
        RECT 112.040 94.275 112.880 94.535 ;
        RECT 117.680 99.000 118.520 99.720 ;
        RECT 124.200 99.490 124.550 101.650 ;
        RECT 113.920 94.275 114.760 94.535 ;
        RECT 124.200 94.990 124.550 97.150 ;
        RECT 40.300 93.000 41.140 93.260 ;
        RECT 42.180 93.000 43.020 93.260 ;
        RECT 47.820 93.040 48.660 93.300 ;
        RECT 49.700 93.040 50.540 93.300 ;
        RECT 51.580 93.040 52.420 93.300 ;
        RECT 40.300 89.950 41.140 90.660 ;
        RECT 42.180 89.950 43.020 90.660 ;
        RECT 37.430 88.510 37.700 89.510 ;
        RECT 39.860 87.800 40.370 88.320 ;
        RECT 34.880 85.640 35.800 86.560 ;
        RECT 44.060 89.950 44.900 90.660 ;
        RECT 38.630 85.640 39.550 86.560 ;
        RECT 39.860 86.050 40.370 86.570 ;
        RECT 40.300 81.665 41.140 82.375 ;
        RECT 41.440 81.230 41.910 82.810 ;
        RECT 43.670 87.820 44.180 88.330 ;
        RECT 45.225 89.610 45.625 91.010 ;
        RECT 45.940 89.950 46.780 90.660 ;
        RECT 47.820 89.950 48.660 90.660 ;
        RECT 62.960 93.000 63.800 93.260 ;
        RECT 64.840 93.000 65.680 93.260 ;
        RECT 70.480 93.040 71.320 93.300 ;
        RECT 72.360 93.040 73.200 93.300 ;
        RECT 74.240 93.040 75.080 93.300 ;
        RECT 49.700 89.950 50.540 90.660 ;
        RECT 48.640 87.820 49.140 88.320 ;
        RECT 51.580 89.950 52.420 90.660 ;
        RECT 53.460 90.040 54.010 90.490 ;
        RECT 55.040 90.130 55.300 90.390 ;
        RECT 56.220 89.940 56.570 92.100 ;
        RECT 62.960 89.950 63.800 90.660 ;
        RECT 64.840 89.950 65.680 90.660 ;
        RECT 50.520 87.820 51.020 88.320 ;
        RECT 43.670 86.040 44.180 86.560 ;
        RECT 42.180 81.665 43.020 82.375 ;
        RECT 48.640 86.120 49.140 86.620 ;
        RECT 50.520 86.120 51.020 86.620 ;
        RECT 56.220 85.440 56.570 87.600 ;
        RECT 59.490 88.510 59.760 89.510 ;
        RECT 62.520 87.800 63.030 88.320 ;
        RECT 57.540 85.640 58.460 86.560 ;
        RECT 66.720 89.950 67.560 90.660 ;
        RECT 61.290 85.640 62.210 86.560 ;
        RECT 62.520 86.050 63.030 86.570 ;
        RECT 44.060 81.665 44.900 82.375 ;
        RECT 45.940 81.665 46.780 82.375 ;
        RECT 47.820 81.660 48.660 82.380 ;
        RECT 44.060 76.935 44.900 77.195 ;
        RECT 49.700 81.660 50.540 82.380 ;
        RECT 56.220 82.150 56.570 84.310 ;
        RECT 62.960 81.665 63.800 82.375 ;
        RECT 45.940 76.935 46.780 77.195 ;
        RECT 56.220 77.650 56.570 79.810 ;
        RECT 64.100 81.230 64.570 82.810 ;
        RECT 66.330 87.820 66.840 88.330 ;
        RECT 67.885 89.610 68.285 91.010 ;
        RECT 68.600 89.950 69.440 90.660 ;
        RECT 70.480 89.950 71.320 90.660 ;
        RECT 85.620 93.000 86.460 93.260 ;
        RECT 87.500 93.000 88.340 93.260 ;
        RECT 93.140 93.040 93.980 93.300 ;
        RECT 95.020 93.040 95.860 93.300 ;
        RECT 96.900 93.040 97.740 93.300 ;
        RECT 72.360 89.950 73.200 90.660 ;
        RECT 71.300 87.820 71.800 88.320 ;
        RECT 74.240 89.950 75.080 90.660 ;
        RECT 76.120 90.040 76.670 90.490 ;
        RECT 77.700 90.130 77.960 90.390 ;
        RECT 78.880 89.940 79.230 92.100 ;
        RECT 85.620 89.950 86.460 90.660 ;
        RECT 87.500 89.950 88.340 90.660 ;
        RECT 73.180 87.820 73.680 88.320 ;
        RECT 66.330 86.040 66.840 86.560 ;
        RECT 64.840 81.665 65.680 82.375 ;
        RECT 71.300 86.120 71.800 86.620 ;
        RECT 73.180 86.120 73.680 86.620 ;
        RECT 78.880 85.440 79.230 87.600 ;
        RECT 82.750 88.510 83.020 89.510 ;
        RECT 85.180 87.800 85.690 88.320 ;
        RECT 80.200 85.640 81.120 86.560 ;
        RECT 89.380 89.950 90.220 90.660 ;
        RECT 83.950 85.640 84.870 86.560 ;
        RECT 85.180 86.050 85.690 86.570 ;
        RECT 66.720 81.665 67.560 82.375 ;
        RECT 68.600 81.665 69.440 82.375 ;
        RECT 70.480 81.660 71.320 82.380 ;
        RECT 66.720 76.935 67.560 77.195 ;
        RECT 72.360 81.660 73.200 82.380 ;
        RECT 78.880 82.150 79.230 84.310 ;
        RECT 85.620 81.665 86.460 82.375 ;
        RECT 68.600 76.935 69.440 77.195 ;
        RECT 78.880 77.650 79.230 79.810 ;
        RECT 86.760 81.230 87.230 82.810 ;
        RECT 88.990 87.820 89.500 88.330 ;
        RECT 90.545 89.610 90.945 91.010 ;
        RECT 91.260 89.950 92.100 90.660 ;
        RECT 93.140 89.950 93.980 90.660 ;
        RECT 108.280 93.000 109.120 93.260 ;
        RECT 110.160 93.000 111.000 93.260 ;
        RECT 115.800 93.040 116.640 93.300 ;
        RECT 117.680 93.040 118.520 93.300 ;
        RECT 119.560 93.040 120.400 93.300 ;
        RECT 95.020 89.950 95.860 90.660 ;
        RECT 93.960 87.820 94.460 88.320 ;
        RECT 96.900 89.950 97.740 90.660 ;
        RECT 98.780 90.040 99.330 90.490 ;
        RECT 100.360 90.130 100.620 90.390 ;
        RECT 101.540 89.940 101.890 92.100 ;
        RECT 108.280 89.950 109.120 90.660 ;
        RECT 110.160 89.950 111.000 90.660 ;
        RECT 95.840 87.820 96.340 88.320 ;
        RECT 88.990 86.040 89.500 86.560 ;
        RECT 87.500 81.665 88.340 82.375 ;
        RECT 93.960 86.120 94.460 86.620 ;
        RECT 95.840 86.120 96.340 86.620 ;
        RECT 101.540 85.440 101.890 87.600 ;
        RECT 104.810 88.510 105.080 89.510 ;
        RECT 107.840 87.800 108.350 88.320 ;
        RECT 102.860 85.640 103.780 86.560 ;
        RECT 112.040 89.950 112.880 90.660 ;
        RECT 106.610 85.640 107.530 86.560 ;
        RECT 107.840 86.050 108.350 86.570 ;
        RECT 89.380 81.665 90.220 82.375 ;
        RECT 91.260 81.665 92.100 82.375 ;
        RECT 93.140 81.660 93.980 82.380 ;
        RECT 89.380 76.935 90.220 77.195 ;
        RECT 95.020 81.660 95.860 82.380 ;
        RECT 101.540 82.150 101.890 84.310 ;
        RECT 108.280 81.665 109.120 82.375 ;
        RECT 91.260 76.935 92.100 77.195 ;
        RECT 101.540 77.650 101.890 79.810 ;
        RECT 109.420 81.230 109.890 82.810 ;
        RECT 111.650 87.820 112.160 88.330 ;
        RECT 113.205 89.610 113.605 91.010 ;
        RECT 113.920 89.950 114.760 90.660 ;
        RECT 115.800 89.950 116.640 90.660 ;
        RECT 117.680 89.950 118.520 90.660 ;
        RECT 116.620 87.820 117.120 88.320 ;
        RECT 119.560 89.950 120.400 90.660 ;
        RECT 121.440 90.040 121.990 90.490 ;
        RECT 123.020 90.130 123.280 90.390 ;
        RECT 124.200 89.940 124.550 92.100 ;
        RECT 118.500 87.820 119.000 88.320 ;
        RECT 111.650 86.040 112.160 86.560 ;
        RECT 110.160 81.665 111.000 82.375 ;
        RECT 116.620 86.120 117.120 86.620 ;
        RECT 118.500 86.120 119.000 86.620 ;
        RECT 124.200 85.440 124.550 87.600 ;
        RECT 112.040 81.665 112.880 82.375 ;
        RECT 113.920 81.665 114.760 82.375 ;
        RECT 115.800 81.660 116.640 82.380 ;
        RECT 112.040 76.935 112.880 77.195 ;
        RECT 117.680 81.660 118.520 82.380 ;
        RECT 124.200 82.150 124.550 84.310 ;
        RECT 113.920 76.935 114.760 77.195 ;
        RECT 124.200 77.650 124.550 79.810 ;
        RECT 40.300 75.660 41.140 75.920 ;
        RECT 42.180 75.660 43.020 75.920 ;
        RECT 47.820 75.700 48.660 75.960 ;
        RECT 49.700 75.700 50.540 75.960 ;
        RECT 51.580 75.700 52.420 75.960 ;
        RECT 40.300 72.610 41.140 73.320 ;
        RECT 42.180 72.610 43.020 73.320 ;
        RECT 38.030 71.170 38.300 72.170 ;
        RECT 39.860 70.460 40.370 70.980 ;
        RECT 34.880 68.300 35.800 69.220 ;
        RECT 44.060 72.610 44.900 73.320 ;
        RECT 38.630 68.300 39.550 69.220 ;
        RECT 39.860 68.710 40.370 69.230 ;
        RECT 40.300 64.325 41.140 65.035 ;
        RECT 41.440 63.890 41.910 65.470 ;
        RECT 43.670 70.480 44.180 70.990 ;
        RECT 45.225 72.270 45.625 73.670 ;
        RECT 45.940 72.610 46.780 73.320 ;
        RECT 47.820 72.610 48.660 73.320 ;
        RECT 62.960 75.660 63.800 75.920 ;
        RECT 64.840 75.660 65.680 75.920 ;
        RECT 70.480 75.700 71.320 75.960 ;
        RECT 72.360 75.700 73.200 75.960 ;
        RECT 74.240 75.700 75.080 75.960 ;
        RECT 49.700 72.610 50.540 73.320 ;
        RECT 48.640 70.480 49.140 70.980 ;
        RECT 51.580 72.610 52.420 73.320 ;
        RECT 53.460 72.700 54.010 73.150 ;
        RECT 55.040 72.790 55.300 73.050 ;
        RECT 56.220 72.600 56.570 74.760 ;
        RECT 62.960 72.610 63.800 73.320 ;
        RECT 64.840 72.610 65.680 73.320 ;
        RECT 50.520 70.480 51.020 70.980 ;
        RECT 43.670 68.700 44.180 69.220 ;
        RECT 42.180 64.325 43.020 65.035 ;
        RECT 48.640 68.780 49.140 69.280 ;
        RECT 50.520 68.780 51.020 69.280 ;
        RECT 56.220 68.100 56.570 70.260 ;
        RECT 58.890 71.170 59.160 72.170 ;
        RECT 62.520 70.460 63.030 70.980 ;
        RECT 57.540 68.300 58.460 69.220 ;
        RECT 66.720 72.610 67.560 73.320 ;
        RECT 61.290 68.300 62.210 69.220 ;
        RECT 62.520 68.710 63.030 69.230 ;
        RECT 44.060 64.325 44.900 65.035 ;
        RECT 45.940 64.325 46.780 65.035 ;
        RECT 47.820 64.320 48.660 65.040 ;
        RECT 44.060 59.595 44.900 59.855 ;
        RECT 49.700 64.320 50.540 65.040 ;
        RECT 56.220 64.810 56.570 66.970 ;
        RECT 62.960 64.325 63.800 65.035 ;
        RECT 45.940 59.595 46.780 59.855 ;
        RECT 56.220 60.310 56.570 62.470 ;
        RECT 64.100 63.890 64.570 65.470 ;
        RECT 66.330 70.480 66.840 70.990 ;
        RECT 67.885 72.270 68.285 73.670 ;
        RECT 68.600 72.610 69.440 73.320 ;
        RECT 70.480 72.610 71.320 73.320 ;
        RECT 85.620 75.660 86.460 75.920 ;
        RECT 87.500 75.660 88.340 75.920 ;
        RECT 93.140 75.700 93.980 75.960 ;
        RECT 95.020 75.700 95.860 75.960 ;
        RECT 96.900 75.700 97.740 75.960 ;
        RECT 72.360 72.610 73.200 73.320 ;
        RECT 71.300 70.480 71.800 70.980 ;
        RECT 74.240 72.610 75.080 73.320 ;
        RECT 76.120 72.700 76.670 73.150 ;
        RECT 77.700 72.790 77.960 73.050 ;
        RECT 78.880 72.600 79.230 74.760 ;
        RECT 85.620 72.610 86.460 73.320 ;
        RECT 87.500 72.610 88.340 73.320 ;
        RECT 73.180 70.480 73.680 70.980 ;
        RECT 66.330 68.700 66.840 69.220 ;
        RECT 64.840 64.325 65.680 65.035 ;
        RECT 71.300 68.780 71.800 69.280 ;
        RECT 73.180 68.780 73.680 69.280 ;
        RECT 78.880 68.100 79.230 70.260 ;
        RECT 83.350 71.170 83.620 72.170 ;
        RECT 85.180 70.460 85.690 70.980 ;
        RECT 80.200 68.300 81.120 69.220 ;
        RECT 89.380 72.610 90.220 73.320 ;
        RECT 83.950 68.300 84.870 69.220 ;
        RECT 85.180 68.710 85.690 69.230 ;
        RECT 66.720 64.325 67.560 65.035 ;
        RECT 68.600 64.325 69.440 65.035 ;
        RECT 70.480 64.320 71.320 65.040 ;
        RECT 66.720 59.595 67.560 59.855 ;
        RECT 72.360 64.320 73.200 65.040 ;
        RECT 78.880 64.810 79.230 66.970 ;
        RECT 85.620 64.325 86.460 65.035 ;
        RECT 68.600 59.595 69.440 59.855 ;
        RECT 78.880 60.310 79.230 62.470 ;
        RECT 86.760 63.890 87.230 65.470 ;
        RECT 88.990 70.480 89.500 70.990 ;
        RECT 90.545 72.270 90.945 73.670 ;
        RECT 91.260 72.610 92.100 73.320 ;
        RECT 93.140 72.610 93.980 73.320 ;
        RECT 108.280 75.660 109.120 75.920 ;
        RECT 110.160 75.660 111.000 75.920 ;
        RECT 115.800 75.700 116.640 75.960 ;
        RECT 117.680 75.700 118.520 75.960 ;
        RECT 119.560 75.700 120.400 75.960 ;
        RECT 95.020 72.610 95.860 73.320 ;
        RECT 93.960 70.480 94.460 70.980 ;
        RECT 96.900 72.610 97.740 73.320 ;
        RECT 98.780 72.700 99.330 73.150 ;
        RECT 100.360 72.790 100.620 73.050 ;
        RECT 101.540 72.600 101.890 74.760 ;
        RECT 108.280 72.610 109.120 73.320 ;
        RECT 110.160 72.610 111.000 73.320 ;
        RECT 95.840 70.480 96.340 70.980 ;
        RECT 88.990 68.700 89.500 69.220 ;
        RECT 87.500 64.325 88.340 65.035 ;
        RECT 93.960 68.780 94.460 69.280 ;
        RECT 95.840 68.780 96.340 69.280 ;
        RECT 101.540 68.100 101.890 70.260 ;
        RECT 104.210 71.170 104.480 72.170 ;
        RECT 107.840 70.460 108.350 70.980 ;
        RECT 102.860 68.300 103.780 69.220 ;
        RECT 112.040 72.610 112.880 73.320 ;
        RECT 106.610 68.300 107.530 69.220 ;
        RECT 107.840 68.710 108.350 69.230 ;
        RECT 89.380 64.325 90.220 65.035 ;
        RECT 91.260 64.325 92.100 65.035 ;
        RECT 93.140 64.320 93.980 65.040 ;
        RECT 89.380 59.595 90.220 59.855 ;
        RECT 95.020 64.320 95.860 65.040 ;
        RECT 101.540 64.810 101.890 66.970 ;
        RECT 108.280 64.325 109.120 65.035 ;
        RECT 91.260 59.595 92.100 59.855 ;
        RECT 101.540 60.310 101.890 62.470 ;
        RECT 109.420 63.890 109.890 65.470 ;
        RECT 111.650 70.480 112.160 70.990 ;
        RECT 113.205 72.270 113.605 73.670 ;
        RECT 113.920 72.610 114.760 73.320 ;
        RECT 115.800 72.610 116.640 73.320 ;
        RECT 117.680 72.610 118.520 73.320 ;
        RECT 116.620 70.480 117.120 70.980 ;
        RECT 119.560 72.610 120.400 73.320 ;
        RECT 121.440 72.700 121.990 73.150 ;
        RECT 123.020 72.790 123.280 73.050 ;
        RECT 124.200 72.600 124.550 74.760 ;
        RECT 118.500 70.480 119.000 70.980 ;
        RECT 111.650 68.700 112.160 69.220 ;
        RECT 110.160 64.325 111.000 65.035 ;
        RECT 116.620 68.780 117.120 69.280 ;
        RECT 118.500 68.780 119.000 69.280 ;
        RECT 124.200 68.100 124.550 70.260 ;
        RECT 112.040 64.325 112.880 65.035 ;
        RECT 113.920 64.325 114.760 65.035 ;
        RECT 115.800 64.320 116.640 65.040 ;
        RECT 112.040 59.595 112.880 59.855 ;
        RECT 117.680 64.320 118.520 65.040 ;
        RECT 124.200 64.810 124.550 66.970 ;
        RECT 113.920 59.595 114.760 59.855 ;
        RECT 124.200 60.310 124.550 62.470 ;
        RECT 56.260 58.620 56.520 58.880 ;
        RECT 78.930 58.620 79.190 58.880 ;
        RECT 101.585 58.620 101.845 58.880 ;
        RECT 124.245 58.620 124.505 58.880 ;
        RECT 40.300 57.660 41.140 57.920 ;
        RECT 42.180 57.660 43.020 57.920 ;
        RECT 47.820 57.700 48.660 57.960 ;
        RECT 49.700 57.700 50.540 57.960 ;
        RECT 51.580 57.700 52.420 57.960 ;
        RECT 40.300 54.610 41.140 55.320 ;
        RECT 42.180 54.610 43.020 55.320 ;
        RECT 39.860 52.460 40.370 52.980 ;
        RECT 44.060 54.610 44.900 55.320 ;
        RECT 39.860 50.710 40.370 51.230 ;
        RECT 40.300 46.325 41.140 47.035 ;
        RECT 41.440 45.890 41.910 47.470 ;
        RECT 43.670 52.480 44.180 52.990 ;
        RECT 45.225 54.270 45.625 55.670 ;
        RECT 47.820 54.610 48.660 55.320 ;
        RECT 62.960 57.660 63.800 57.920 ;
        RECT 64.840 57.660 65.680 57.920 ;
        RECT 70.480 57.700 71.320 57.960 ;
        RECT 72.360 57.700 73.200 57.960 ;
        RECT 74.240 57.700 75.080 57.960 ;
        RECT 49.700 54.610 50.540 55.320 ;
        RECT 48.640 52.480 49.140 52.980 ;
        RECT 51.580 54.610 52.420 55.320 ;
        RECT 62.960 54.610 63.800 55.320 ;
        RECT 64.840 54.610 65.680 55.320 ;
        RECT 50.520 52.480 51.020 52.980 ;
        RECT 62.520 52.460 63.030 52.980 ;
        RECT 43.670 50.700 44.180 51.220 ;
        RECT 48.640 50.780 49.140 51.280 ;
        RECT 50.520 50.780 51.020 51.280 ;
        RECT 66.720 54.610 67.560 55.320 ;
        RECT 62.520 50.710 63.030 51.230 ;
        RECT 44.060 46.325 44.900 47.035 ;
        RECT 45.940 46.325 46.780 47.035 ;
        RECT 47.820 46.320 48.660 47.040 ;
        RECT 44.060 41.595 44.900 41.855 ;
        RECT 49.700 46.320 50.540 47.040 ;
        RECT 62.960 46.325 63.800 47.035 ;
        RECT 45.940 41.595 46.780 41.855 ;
        RECT 64.100 45.890 64.570 47.470 ;
        RECT 66.330 52.480 66.840 52.990 ;
        RECT 67.885 54.270 68.285 55.670 ;
        RECT 70.480 54.610 71.320 55.320 ;
        RECT 85.620 57.660 86.460 57.920 ;
        RECT 87.500 57.660 88.340 57.920 ;
        RECT 93.140 57.700 93.980 57.960 ;
        RECT 95.020 57.700 95.860 57.960 ;
        RECT 96.900 57.700 97.740 57.960 ;
        RECT 72.360 54.610 73.200 55.320 ;
        RECT 71.300 52.480 71.800 52.980 ;
        RECT 74.240 54.610 75.080 55.320 ;
        RECT 85.620 54.610 86.460 55.320 ;
        RECT 87.500 54.610 88.340 55.320 ;
        RECT 73.180 52.480 73.680 52.980 ;
        RECT 85.180 52.460 85.690 52.980 ;
        RECT 66.330 50.700 66.840 51.220 ;
        RECT 71.300 50.780 71.800 51.280 ;
        RECT 73.180 50.780 73.680 51.280 ;
        RECT 89.380 54.610 90.220 55.320 ;
        RECT 85.180 50.710 85.690 51.230 ;
        RECT 66.720 46.325 67.560 47.035 ;
        RECT 68.600 46.325 69.440 47.035 ;
        RECT 70.480 46.320 71.320 47.040 ;
        RECT 66.720 41.595 67.560 41.855 ;
        RECT 72.360 46.320 73.200 47.040 ;
        RECT 85.620 46.325 86.460 47.035 ;
        RECT 68.600 41.595 69.440 41.855 ;
        RECT 86.760 45.890 87.230 47.470 ;
        RECT 88.990 52.480 89.500 52.990 ;
        RECT 90.545 54.270 90.945 55.670 ;
        RECT 93.140 54.610 93.980 55.320 ;
        RECT 108.280 57.660 109.120 57.920 ;
        RECT 110.160 57.660 111.000 57.920 ;
        RECT 115.800 57.700 116.640 57.960 ;
        RECT 117.680 57.700 118.520 57.960 ;
        RECT 119.560 57.700 120.400 57.960 ;
        RECT 95.020 54.610 95.860 55.320 ;
        RECT 93.960 52.480 94.460 52.980 ;
        RECT 96.900 54.610 97.740 55.320 ;
        RECT 108.280 54.610 109.120 55.320 ;
        RECT 110.160 54.610 111.000 55.320 ;
        RECT 95.840 52.480 96.340 52.980 ;
        RECT 107.840 52.460 108.350 52.980 ;
        RECT 88.990 50.700 89.500 51.220 ;
        RECT 93.960 50.780 94.460 51.280 ;
        RECT 95.840 50.780 96.340 51.280 ;
        RECT 112.040 54.610 112.880 55.320 ;
        RECT 107.840 50.710 108.350 51.230 ;
        RECT 89.380 46.325 90.220 47.035 ;
        RECT 91.260 46.325 92.100 47.035 ;
        RECT 93.140 46.320 93.980 47.040 ;
        RECT 89.380 41.595 90.220 41.855 ;
        RECT 95.020 46.320 95.860 47.040 ;
        RECT 108.280 46.325 109.120 47.035 ;
        RECT 91.260 41.595 92.100 41.855 ;
        RECT 109.420 45.890 109.890 47.470 ;
        RECT 111.650 52.480 112.160 52.990 ;
        RECT 113.205 54.270 113.605 55.670 ;
        RECT 115.800 54.610 116.640 55.320 ;
        RECT 117.680 54.610 118.520 55.320 ;
        RECT 116.620 52.480 117.120 52.980 ;
        RECT 119.560 54.610 120.400 55.320 ;
        RECT 118.500 52.480 119.000 52.980 ;
        RECT 111.650 50.700 112.160 51.220 ;
        RECT 116.620 50.780 117.120 51.280 ;
        RECT 118.500 50.780 119.000 51.280 ;
        RECT 112.040 46.325 112.880 47.035 ;
        RECT 113.920 46.325 114.760 47.035 ;
        RECT 115.800 46.320 116.640 47.040 ;
        RECT 112.040 41.595 112.880 41.855 ;
        RECT 117.680 46.320 118.520 47.040 ;
        RECT 113.920 41.595 114.760 41.855 ;
      LAYER met2 ;
        RECT 76.380 187.620 76.640 187.940 ;
        RECT 93.400 187.620 93.660 187.940 ;
        RECT 74.540 187.280 74.800 187.600 ;
        RECT 57.060 184.900 57.320 185.220 ;
        RECT 58.440 184.900 58.700 185.220 ;
        RECT 62.580 184.900 62.840 185.220 ;
        RECT 65.800 184.900 66.060 185.220 ;
        RECT 69.940 184.900 70.200 185.220 ;
        RECT 73.160 184.900 73.420 185.220 ;
        RECT 55.220 182.860 55.480 183.180 ;
        RECT 54.300 181.840 54.560 182.160 ;
        RECT 53.840 181.500 54.100 181.820 ;
        RECT 52.460 179.120 52.720 179.440 ;
        RECT 49.700 178.780 49.960 179.100 ;
        RECT 49.760 178.080 49.900 178.780 ;
        RECT 49.700 177.760 49.960 178.080 ;
        RECT 51.540 176.915 51.800 177.060 ;
        RECT 51.530 176.800 51.810 176.915 ;
        RECT 51.530 176.660 52.200 176.800 ;
        RECT 51.530 176.545 51.810 176.660 ;
        RECT 52.060 174.340 52.200 176.660 ;
        RECT 52.520 174.680 52.660 179.120 ;
        RECT 53.900 179.100 54.040 181.500 ;
        RECT 54.360 179.780 54.500 181.840 ;
        RECT 54.300 179.460 54.560 179.780 ;
        RECT 53.840 178.780 54.100 179.100 ;
        RECT 52.460 174.360 52.720 174.680 ;
        RECT 52.000 174.020 52.260 174.340 ;
        RECT 44.640 171.640 44.900 171.960 ;
        RECT 44.700 159.040 44.840 171.640 ;
        RECT 53.900 166.180 54.040 178.780 ;
        RECT 55.280 174.340 55.420 182.860 ;
        RECT 56.600 182.520 56.860 182.840 ;
        RECT 56.660 176.720 56.800 182.520 ;
        RECT 56.600 176.400 56.860 176.720 ;
        RECT 55.220 174.020 55.480 174.340 ;
        RECT 56.140 173.340 56.400 173.660 ;
        RECT 54.300 171.300 54.560 171.620 ;
        RECT 54.360 167.200 54.500 171.300 ;
        RECT 54.760 170.620 55.020 170.940 ;
        RECT 54.820 167.200 54.960 170.620 ;
        RECT 55.220 168.580 55.480 168.900 ;
        RECT 54.300 166.880 54.560 167.200 ;
        RECT 54.760 166.880 55.020 167.200 ;
        RECT 54.820 166.520 54.960 166.880 ;
        RECT 55.280 166.520 55.420 168.580 ;
        RECT 54.760 166.200 55.020 166.520 ;
        RECT 55.220 166.200 55.480 166.520 ;
        RECT 53.840 165.860 54.100 166.180 ;
        RECT 53.900 163.120 54.040 165.860 ;
        RECT 53.840 162.800 54.100 163.120 ;
        RECT 54.820 161.760 54.960 166.200 ;
        RECT 55.280 163.800 55.420 166.200 ;
        RECT 55.220 163.480 55.480 163.800 ;
        RECT 55.220 162.460 55.480 162.780 ;
        RECT 54.760 161.440 55.020 161.760 ;
        RECT 52.920 160.760 53.180 161.080 ;
        RECT 44.640 158.720 44.900 159.040 ;
        RECT 52.980 158.360 53.120 160.760 ;
        RECT 55.280 160.740 55.420 162.460 ;
        RECT 55.220 160.420 55.480 160.740 ;
        RECT 56.200 159.040 56.340 173.340 ;
        RECT 57.120 172.640 57.260 184.900 ;
        RECT 57.520 179.460 57.780 179.780 ;
        RECT 57.580 177.060 57.720 179.460 ;
        RECT 58.500 178.080 58.640 184.900 ;
        RECT 62.120 182.520 62.380 182.840 ;
        RECT 60.280 179.350 60.540 179.440 ;
        RECT 61.200 179.350 61.460 179.440 ;
        RECT 60.280 179.210 61.460 179.350 ;
        RECT 60.280 179.120 60.540 179.210 ;
        RECT 61.200 179.120 61.460 179.210 ;
        RECT 62.180 178.080 62.320 182.520 ;
        RECT 62.640 180.800 62.780 184.900 ;
        RECT 63.960 184.560 64.220 184.880 ;
        RECT 63.500 182.180 63.760 182.500 ;
        RECT 62.580 180.480 62.840 180.800 ;
        RECT 62.580 179.460 62.840 179.780 ;
        RECT 58.440 177.760 58.700 178.080 ;
        RECT 62.120 177.760 62.380 178.080 ;
        RECT 57.520 176.740 57.780 177.060 ;
        RECT 60.740 176.740 61.000 177.060 ;
        RECT 61.200 176.740 61.460 177.060 ;
        RECT 57.060 172.320 57.320 172.640 ;
        RECT 57.580 165.840 57.720 176.740 ;
        RECT 60.800 175.360 60.940 176.740 ;
        RECT 60.740 175.040 61.000 175.360 ;
        RECT 61.260 174.680 61.400 176.740 ;
        RECT 62.180 176.120 62.320 177.760 ;
        RECT 61.720 175.980 62.320 176.120 ;
        RECT 61.200 174.360 61.460 174.680 ;
        RECT 58.900 174.020 59.160 174.340 ;
        RECT 59.360 174.195 59.620 174.340 ;
        RECT 58.440 173.340 58.700 173.660 ;
        RECT 57.980 167.900 58.240 168.220 ;
        RECT 57.520 165.520 57.780 165.840 ;
        RECT 57.580 165.355 57.720 165.520 ;
        RECT 57.510 164.985 57.790 165.355 ;
        RECT 58.040 161.760 58.180 167.900 ;
        RECT 58.500 166.180 58.640 173.340 ;
        RECT 58.960 171.960 59.100 174.020 ;
        RECT 59.350 173.825 59.630 174.195 ;
        RECT 58.900 171.640 59.160 171.960 ;
        RECT 60.740 171.530 61.000 171.620 ;
        RECT 61.260 171.530 61.400 174.360 ;
        RECT 60.740 171.390 61.400 171.530 ;
        RECT 60.740 171.300 61.000 171.390 ;
        RECT 60.800 169.240 60.940 171.300 ;
        RECT 60.740 168.920 61.000 169.240 ;
        RECT 58.440 165.860 58.700 166.180 ;
        RECT 59.820 165.860 60.080 166.180 ;
        RECT 59.880 165.500 60.020 165.860 ;
        RECT 59.820 165.180 60.080 165.500 ;
        RECT 59.880 163.460 60.020 165.180 ;
        RECT 59.820 163.140 60.080 163.460 ;
        RECT 57.980 161.440 58.240 161.760 ;
        RECT 61.720 159.040 61.860 175.980 ;
        RECT 56.140 158.720 56.400 159.040 ;
        RECT 61.660 158.720 61.920 159.040 ;
        RECT 62.640 158.700 62.780 179.460 ;
        RECT 63.560 178.080 63.700 182.180 ;
        RECT 63.500 177.760 63.760 178.080 ;
        RECT 63.560 176.380 63.700 177.760 ;
        RECT 63.500 176.060 63.760 176.380 ;
        RECT 63.500 173.340 63.760 173.660 ;
        RECT 63.560 164.480 63.700 173.340 ;
        RECT 64.020 169.920 64.160 184.560 ;
        RECT 64.880 180.480 65.140 180.800 ;
        RECT 64.940 179.780 65.080 180.480 ;
        RECT 64.880 179.460 65.140 179.780 ;
        RECT 65.340 178.780 65.600 179.100 ;
        RECT 65.400 177.740 65.540 178.780 ;
        RECT 65.340 177.420 65.600 177.740 ;
        RECT 65.860 173.660 66.000 184.900 ;
        RECT 67.180 183.200 67.440 183.520 ;
        RECT 67.240 180.120 67.380 183.200 ;
        RECT 70.000 182.240 70.140 184.900 ;
        RECT 73.220 183.520 73.360 184.900 ;
        RECT 73.620 184.560 73.880 184.880 ;
        RECT 73.160 183.200 73.420 183.520 ;
        RECT 70.000 182.100 70.600 182.240 ;
        RECT 72.700 182.180 72.960 182.500 ;
        RECT 66.260 179.800 66.520 180.120 ;
        RECT 67.180 179.800 67.440 180.120 ;
        RECT 66.320 177.060 66.460 179.800 ;
        RECT 66.720 178.780 66.980 179.100 ;
        RECT 66.260 176.740 66.520 177.060 ;
        RECT 65.800 173.340 66.060 173.660 ;
        RECT 66.260 173.340 66.520 173.660 ;
        RECT 64.420 171.980 64.680 172.300 ;
        RECT 63.960 169.600 64.220 169.920 ;
        RECT 64.480 168.560 64.620 171.980 ;
        RECT 66.320 171.960 66.460 173.340 ;
        RECT 65.800 171.640 66.060 171.960 ;
        RECT 66.260 171.640 66.520 171.960 ;
        RECT 64.420 168.240 64.680 168.560 ;
        RECT 63.500 164.160 63.760 164.480 ;
        RECT 64.480 159.040 64.620 168.240 ;
        RECT 65.860 167.820 66.000 171.640 ;
        RECT 66.780 171.620 66.920 178.780 ;
        RECT 67.640 174.020 67.900 174.340 ;
        RECT 69.940 174.020 70.200 174.340 ;
        RECT 66.720 171.300 66.980 171.620 ;
        RECT 67.700 169.240 67.840 174.020 ;
        RECT 68.100 173.340 68.360 173.660 ;
        RECT 68.160 172.640 68.300 173.340 ;
        RECT 68.100 172.320 68.360 172.640 ;
        RECT 70.000 172.300 70.140 174.020 ;
        RECT 69.940 171.980 70.200 172.300 ;
        RECT 68.100 170.620 68.360 170.940 ;
        RECT 67.640 168.920 67.900 169.240 ;
        RECT 68.160 168.900 68.300 170.620 ;
        RECT 68.100 168.580 68.360 168.900 ;
        RECT 68.560 168.580 68.820 168.900 ;
        RECT 68.620 167.820 68.760 168.580 ;
        RECT 65.860 167.680 68.760 167.820 ;
        RECT 65.860 163.460 66.000 167.680 ;
        RECT 68.620 167.200 68.760 167.680 ;
        RECT 68.560 166.880 68.820 167.200 ;
        RECT 67.170 164.985 67.450 165.355 ;
        RECT 67.240 164.140 67.380 164.985 ;
        RECT 67.180 163.820 67.440 164.140 ;
        RECT 69.480 163.480 69.740 163.800 ;
        RECT 65.340 163.140 65.600 163.460 ;
        RECT 65.800 163.140 66.060 163.460 ;
        RECT 65.400 162.780 65.540 163.140 ;
        RECT 65.340 162.460 65.600 162.780 ;
        RECT 65.400 161.760 65.540 162.460 ;
        RECT 65.340 161.440 65.600 161.760 ;
        RECT 65.860 161.420 66.000 163.140 ;
        RECT 65.800 161.100 66.060 161.420 ;
        RECT 69.540 161.080 69.680 163.480 ;
        RECT 69.940 163.140 70.200 163.460 ;
        RECT 69.480 160.760 69.740 161.080 ;
        RECT 70.000 160.740 70.140 163.140 ;
        RECT 70.460 161.760 70.600 182.100 ;
        RECT 72.760 181.820 72.900 182.180 ;
        RECT 72.700 181.500 72.960 181.820 ;
        RECT 70.850 177.225 71.130 177.595 ;
        RECT 70.920 164.140 71.060 177.225 ;
        RECT 72.760 175.020 72.900 181.500 ;
        RECT 73.160 177.080 73.420 177.400 ;
        RECT 72.700 174.700 72.960 175.020 ;
        RECT 72.240 174.020 72.500 174.340 ;
        RECT 72.300 172.640 72.440 174.020 ;
        RECT 72.240 172.320 72.500 172.640 ;
        RECT 72.700 171.980 72.960 172.300 ;
        RECT 73.220 172.155 73.360 177.080 ;
        RECT 72.760 169.240 72.900 171.980 ;
        RECT 73.150 171.785 73.430 172.155 ;
        RECT 72.700 168.920 72.960 169.240 ;
        RECT 71.780 167.900 72.040 168.220 ;
        RECT 71.840 166.860 71.980 167.900 ;
        RECT 71.780 166.540 72.040 166.860 ;
        RECT 72.700 165.180 72.960 165.500 ;
        RECT 70.860 163.820 71.120 164.140 ;
        RECT 72.760 163.460 72.900 165.180 ;
        RECT 73.150 163.625 73.430 163.995 ;
        RECT 73.160 163.480 73.420 163.625 ;
        RECT 72.700 163.140 72.960 163.460 ;
        RECT 73.680 161.760 73.820 184.560 ;
        RECT 74.600 183.520 74.740 187.280 ;
        RECT 75.920 184.900 76.180 185.220 ;
        RECT 74.540 183.200 74.800 183.520 ;
        RECT 75.000 183.200 75.260 183.520 ;
        RECT 75.060 178.840 75.200 183.200 ;
        RECT 75.460 179.120 75.720 179.440 ;
        RECT 74.600 178.700 75.200 178.840 ;
        RECT 74.600 176.970 74.740 178.700 ;
        RECT 74.600 176.830 75.200 176.970 ;
        RECT 74.080 176.290 74.340 176.380 ;
        RECT 74.080 176.150 74.740 176.290 ;
        RECT 74.080 176.060 74.340 176.150 ;
        RECT 74.080 174.700 74.340 175.020 ;
        RECT 74.140 169.580 74.280 174.700 ;
        RECT 74.080 169.260 74.340 169.580 ;
        RECT 74.600 167.820 74.740 176.150 ;
        RECT 75.060 174.340 75.200 176.830 ;
        RECT 75.000 174.020 75.260 174.340 ;
        RECT 75.060 173.660 75.200 174.020 ;
        RECT 75.000 173.340 75.260 173.660 ;
        RECT 74.140 167.680 74.740 167.820 ;
        RECT 70.400 161.440 70.660 161.760 ;
        RECT 73.620 161.440 73.880 161.760 ;
        RECT 74.140 160.740 74.280 167.680 ;
        RECT 75.520 166.520 75.660 179.120 ;
        RECT 75.980 178.080 76.120 184.900 ;
        RECT 76.440 182.500 76.580 187.620 ;
        RECT 83.740 185.580 84.000 185.900 ;
        RECT 83.280 184.900 83.540 185.220 ;
        RECT 83.340 182.840 83.480 184.900 ;
        RECT 83.800 183.520 83.940 185.580 ;
        RECT 88.800 184.220 89.060 184.540 ;
        RECT 89.260 184.220 89.520 184.540 ;
        RECT 91.100 184.220 91.360 184.540 ;
        RECT 83.740 183.200 84.000 183.520 ;
        RECT 77.300 182.520 77.560 182.840 ;
        RECT 81.900 182.520 82.160 182.840 ;
        RECT 83.280 182.520 83.540 182.840 ;
        RECT 85.580 182.520 85.840 182.840 ;
        RECT 76.380 182.180 76.640 182.500 ;
        RECT 76.840 181.500 77.100 181.820 ;
        RECT 76.900 179.780 77.040 181.500 ;
        RECT 76.840 179.460 77.100 179.780 ;
        RECT 75.920 177.760 76.180 178.080 ;
        RECT 76.380 174.250 76.640 174.340 ;
        RECT 75.980 174.110 76.640 174.250 ;
        RECT 75.980 172.300 76.120 174.110 ;
        RECT 76.380 174.020 76.640 174.110 ;
        RECT 76.380 173.340 76.640 173.660 ;
        RECT 75.920 171.980 76.180 172.300 ;
        RECT 75.980 169.920 76.120 171.980 ;
        RECT 75.920 169.600 76.180 169.920 ;
        RECT 75.460 166.200 75.720 166.520 ;
        RECT 75.000 163.820 75.260 164.140 ;
        RECT 75.060 161.080 75.200 163.820 ;
        RECT 76.440 161.760 76.580 173.340 ;
        RECT 76.840 168.240 77.100 168.560 ;
        RECT 76.380 161.670 76.640 161.760 ;
        RECT 75.980 161.530 76.640 161.670 ;
        RECT 75.000 160.760 75.260 161.080 ;
        RECT 69.940 160.420 70.200 160.740 ;
        RECT 72.240 160.420 72.500 160.740 ;
        RECT 74.080 160.420 74.340 160.740 ;
        RECT 67.640 160.080 67.900 160.400 ;
        RECT 67.180 159.740 67.440 160.060 ;
        RECT 67.240 159.040 67.380 159.740 ;
        RECT 67.700 159.040 67.840 160.080 ;
        RECT 72.300 159.040 72.440 160.420 ;
        RECT 75.060 159.040 75.200 160.760 ;
        RECT 64.420 158.720 64.680 159.040 ;
        RECT 67.180 158.720 67.440 159.040 ;
        RECT 67.640 158.720 67.900 159.040 ;
        RECT 72.240 158.720 72.500 159.040 ;
        RECT 75.000 158.720 75.260 159.040 ;
        RECT 62.580 158.380 62.840 158.700 ;
        RECT 52.920 158.040 53.180 158.360 ;
        RECT 75.980 158.020 76.120 161.530 ;
        RECT 76.380 161.440 76.640 161.530 ;
        RECT 76.900 161.420 77.040 168.240 ;
        RECT 76.840 161.100 77.100 161.420 ;
        RECT 76.380 160.420 76.640 160.740 ;
        RECT 76.440 158.020 76.580 160.420 ;
        RECT 77.360 159.040 77.500 182.520 ;
        RECT 81.960 179.780 82.100 182.520 ;
        RECT 85.640 180.800 85.780 182.520 ;
        RECT 86.040 182.180 86.300 182.500 ;
        RECT 86.500 182.180 86.760 182.500 ;
        RECT 88.860 182.240 89.000 184.220 ;
        RECT 89.320 183.520 89.460 184.220 ;
        RECT 89.260 183.200 89.520 183.520 ;
        RECT 90.640 182.860 90.900 183.180 ;
        RECT 85.580 180.480 85.840 180.800 ;
        RECT 83.280 180.140 83.540 180.460 ;
        RECT 81.900 179.460 82.160 179.780 ;
        RECT 80.060 179.120 80.320 179.440 ;
        RECT 80.120 177.060 80.260 179.120 ;
        RECT 80.060 176.740 80.320 177.060 ;
        RECT 80.980 170.620 81.240 170.940 ;
        RECT 81.440 170.620 81.700 170.940 ;
        RECT 81.040 167.820 81.180 170.620 ;
        RECT 81.500 169.240 81.640 170.620 ;
        RECT 81.440 168.920 81.700 169.240 ;
        RECT 81.440 168.470 81.700 168.560 ;
        RECT 81.960 168.470 82.100 179.460 ;
        RECT 82.360 176.740 82.620 177.060 ;
        RECT 81.440 168.330 82.100 168.470 ;
        RECT 81.440 168.240 81.700 168.330 ;
        RECT 80.580 167.680 81.180 167.820 ;
        RECT 80.580 166.860 80.720 167.680 ;
        RECT 77.760 166.540 78.020 166.860 ;
        RECT 80.520 166.540 80.780 166.860 ;
        RECT 77.820 162.780 77.960 166.540 ;
        RECT 81.440 166.200 81.700 166.520 ;
        RECT 81.500 163.460 81.640 166.200 ;
        RECT 82.420 166.035 82.560 176.740 ;
        RECT 82.810 174.505 83.090 174.875 ;
        RECT 82.820 174.360 83.080 174.505 ;
        RECT 83.340 172.640 83.480 180.140 ;
        RECT 83.740 179.800 84.000 180.120 ;
        RECT 83.280 172.320 83.540 172.640 ;
        RECT 82.820 171.640 83.080 171.960 ;
        RECT 82.880 169.435 83.020 171.640 ;
        RECT 83.340 169.920 83.480 172.320 ;
        RECT 83.280 169.600 83.540 169.920 ;
        RECT 82.810 169.065 83.090 169.435 ;
        RECT 83.800 169.240 83.940 179.800 ;
        RECT 86.100 179.780 86.240 182.180 ;
        RECT 86.560 180.120 86.700 182.180 ;
        RECT 88.860 182.100 89.460 182.240 ;
        RECT 90.180 182.180 90.440 182.500 ;
        RECT 86.500 179.800 86.760 180.120 ;
        RECT 84.660 179.460 84.920 179.780 ;
        RECT 86.040 179.460 86.300 179.780 ;
        RECT 84.200 177.760 84.460 178.080 ;
        RECT 84.260 177.400 84.400 177.760 ;
        RECT 84.720 177.400 84.860 179.460 ;
        RECT 84.200 177.080 84.460 177.400 ;
        RECT 84.660 177.080 84.920 177.400 ;
        RECT 84.260 173.570 84.400 177.080 ;
        RECT 86.100 175.360 86.240 179.460 ;
        RECT 89.320 178.080 89.460 182.100 ;
        RECT 89.720 181.840 89.980 182.160 ;
        RECT 89.780 179.440 89.920 181.840 ;
        RECT 90.240 179.440 90.380 182.180 ;
        RECT 89.720 179.120 89.980 179.440 ;
        RECT 90.180 179.120 90.440 179.440 ;
        RECT 90.700 179.100 90.840 182.860 ;
        RECT 90.640 178.780 90.900 179.100 ;
        RECT 89.260 177.760 89.520 178.080 ;
        RECT 89.250 177.480 89.530 177.595 ;
        RECT 88.860 177.340 89.530 177.480 ;
        RECT 88.860 177.060 89.000 177.340 ;
        RECT 89.250 177.225 89.530 177.340 ;
        RECT 88.800 176.740 89.060 177.060 ;
        RECT 89.260 176.060 89.520 176.380 ;
        RECT 86.040 175.040 86.300 175.360 ;
        RECT 89.320 175.270 89.460 176.060 ;
        RECT 88.860 175.130 89.460 175.270 ;
        RECT 84.660 174.700 84.920 175.020 ;
        RECT 84.720 174.340 84.860 174.700 ;
        RECT 86.030 174.505 86.310 174.875 ;
        RECT 84.660 174.020 84.920 174.340 ;
        RECT 86.100 173.660 86.240 174.505 ;
        RECT 85.120 173.570 85.380 173.660 ;
        RECT 84.260 173.430 85.380 173.570 ;
        RECT 85.120 173.340 85.380 173.430 ;
        RECT 86.040 173.340 86.300 173.660 ;
        RECT 87.880 173.570 88.140 173.660 ;
        RECT 87.480 173.430 88.140 173.570 ;
        RECT 83.740 168.920 84.000 169.240 ;
        RECT 82.820 168.580 83.080 168.900 ;
        RECT 82.350 165.665 82.630 166.035 ;
        RECT 82.420 164.480 82.560 165.665 ;
        RECT 82.360 164.160 82.620 164.480 ;
        RECT 82.880 164.140 83.020 168.580 ;
        RECT 82.820 163.820 83.080 164.140 ;
        RECT 85.180 163.460 85.320 173.340 ;
        RECT 87.480 172.300 87.620 173.430 ;
        RECT 87.880 173.340 88.140 173.430 ;
        RECT 88.340 172.320 88.600 172.640 ;
        RECT 87.420 171.980 87.680 172.300 ;
        RECT 86.960 171.640 87.220 171.960 ;
        RECT 87.020 170.680 87.160 171.640 ;
        RECT 87.410 171.105 87.690 171.475 ;
        RECT 88.400 171.360 88.540 172.320 ;
        RECT 87.940 171.280 88.540 171.360 ;
        RECT 87.880 171.220 88.540 171.280 ;
        RECT 88.860 171.360 89.000 175.130 ;
        RECT 89.720 175.040 89.980 175.360 ;
        RECT 89.260 174.360 89.520 174.680 ;
        RECT 89.320 172.640 89.460 174.360 ;
        RECT 89.260 172.320 89.520 172.640 ;
        RECT 88.860 171.220 89.460 171.360 ;
        RECT 87.480 170.940 87.620 171.105 ;
        RECT 87.880 170.960 88.140 171.220 ;
        RECT 86.560 170.540 87.160 170.680 ;
        RECT 87.420 170.620 87.680 170.940 ;
        RECT 86.560 168.640 86.700 170.540 ;
        RECT 86.950 169.065 87.230 169.435 ;
        RECT 86.960 168.920 87.220 169.065 ;
        RECT 87.880 168.640 88.140 168.900 ;
        RECT 86.560 168.580 88.140 168.640 ;
        RECT 86.560 168.500 88.080 168.580 ;
        RECT 86.560 164.480 86.700 168.500 ;
        RECT 86.500 164.160 86.760 164.480 ;
        RECT 81.440 163.140 81.700 163.460 ;
        RECT 82.360 163.140 82.620 163.460 ;
        RECT 85.120 163.140 85.380 163.460 ;
        RECT 77.760 162.460 78.020 162.780 ;
        RECT 82.420 161.080 82.560 163.140 ;
        RECT 89.320 163.120 89.460 171.220 ;
        RECT 89.780 163.800 89.920 175.040 ;
        RECT 90.180 174.020 90.440 174.340 ;
        RECT 90.240 169.920 90.380 174.020 ;
        RECT 90.180 169.600 90.440 169.920 ;
        RECT 90.180 167.900 90.440 168.220 ;
        RECT 90.240 163.800 90.380 167.900 ;
        RECT 89.720 163.480 89.980 163.800 ;
        RECT 90.180 163.480 90.440 163.800 ;
        RECT 89.260 162.800 89.520 163.120 ;
        RECT 82.360 160.760 82.620 161.080 ;
        RECT 80.980 159.740 81.240 160.060 ;
        RECT 81.440 159.740 81.700 160.060 ;
        RECT 77.300 158.720 77.560 159.040 ;
        RECT 81.040 158.360 81.180 159.740 ;
        RECT 81.500 159.040 81.640 159.740 ;
        RECT 89.320 159.040 89.460 162.800 ;
        RECT 89.720 159.740 89.980 160.060 ;
        RECT 89.780 159.040 89.920 159.740 ;
        RECT 90.700 159.040 90.840 178.780 ;
        RECT 91.160 171.475 91.300 184.220 ;
        RECT 93.460 183.180 93.600 187.620 ;
        RECT 117.320 187.280 117.580 187.600 ;
        RECT 110.420 185.580 110.680 185.900 ;
        RECT 102.140 185.240 102.400 185.560 ;
        RECT 106.740 185.240 107.000 185.560 ;
        RECT 98.460 184.900 98.720 185.220 ;
        RECT 93.860 184.560 94.120 184.880 ;
        RECT 93.920 183.520 94.060 184.560 ;
        RECT 98.520 183.520 98.660 184.900 ;
        RECT 100.760 184.560 101.020 184.880 ;
        RECT 93.860 183.200 94.120 183.520 ;
        RECT 98.460 183.200 98.720 183.520 ;
        RECT 100.300 183.200 100.560 183.520 ;
        RECT 93.400 182.860 93.660 183.180 ;
        RECT 95.700 182.520 95.960 182.840 ;
        RECT 94.780 182.180 95.040 182.500 ;
        RECT 94.840 180.800 94.980 182.180 ;
        RECT 95.240 181.500 95.500 181.820 ;
        RECT 92.020 180.480 92.280 180.800 ;
        RECT 94.780 180.480 95.040 180.800 ;
        RECT 91.560 178.780 91.820 179.100 ;
        RECT 91.090 171.105 91.370 171.475 ;
        RECT 91.620 169.435 91.760 178.780 ;
        RECT 92.080 177.740 92.220 180.480 ;
        RECT 94.320 178.780 94.580 179.100 ;
        RECT 92.020 177.420 92.280 177.740 ;
        RECT 91.550 169.065 91.830 169.435 ;
        RECT 92.080 166.520 92.220 177.420 ;
        RECT 92.940 176.400 93.200 176.720 ;
        RECT 93.000 168.220 93.140 176.400 ;
        RECT 93.400 176.060 93.660 176.380 ;
        RECT 93.460 175.360 93.600 176.060 ;
        RECT 93.400 175.040 93.660 175.360 ;
        RECT 94.380 174.340 94.520 178.780 ;
        RECT 94.320 174.020 94.580 174.340 ;
        RECT 93.860 173.340 94.120 173.660 ;
        RECT 94.320 173.340 94.580 173.660 ;
        RECT 93.920 170.940 94.060 173.340 ;
        RECT 93.860 170.620 94.120 170.940 ;
        RECT 94.380 169.580 94.520 173.340 ;
        RECT 94.840 172.640 94.980 180.480 ;
        RECT 95.300 178.080 95.440 181.500 ;
        RECT 95.240 177.760 95.500 178.080 ;
        RECT 95.240 177.080 95.500 177.400 ;
        RECT 95.300 173.515 95.440 177.080 ;
        RECT 95.230 173.145 95.510 173.515 ;
        RECT 94.780 172.320 95.040 172.640 ;
        RECT 95.300 171.620 95.440 173.145 ;
        RECT 95.240 171.300 95.500 171.620 ;
        RECT 94.780 170.960 95.040 171.280 ;
        RECT 94.320 169.260 94.580 169.580 ;
        RECT 93.400 168.580 93.660 168.900 ;
        RECT 93.860 168.580 94.120 168.900 ;
        RECT 92.940 167.900 93.200 168.220 ;
        RECT 93.460 167.200 93.600 168.580 ;
        RECT 93.400 166.880 93.660 167.200 ;
        RECT 93.920 166.520 94.060 168.580 ;
        RECT 92.020 166.200 92.280 166.520 ;
        RECT 92.480 166.200 92.740 166.520 ;
        RECT 93.860 166.200 94.120 166.520 ;
        RECT 91.560 160.760 91.820 161.080 ;
        RECT 81.440 158.720 81.700 159.040 ;
        RECT 89.260 158.720 89.520 159.040 ;
        RECT 89.720 158.720 89.980 159.040 ;
        RECT 90.640 158.720 90.900 159.040 ;
        RECT 80.980 158.040 81.240 158.360 ;
        RECT 91.620 158.020 91.760 160.760 ;
        RECT 92.080 160.740 92.220 166.200 ;
        RECT 92.540 164.480 92.680 166.200 ;
        RECT 92.480 164.160 92.740 164.480 ;
        RECT 94.840 163.800 94.980 170.960 ;
        RECT 94.780 163.480 95.040 163.800 ;
        RECT 95.300 163.460 95.440 171.300 ;
        RECT 95.760 169.240 95.900 182.520 ;
        RECT 98.920 182.180 99.180 182.500 ;
        RECT 96.160 179.460 96.420 179.780 ;
        RECT 96.220 177.740 96.360 179.460 ;
        RECT 96.620 177.760 96.880 178.080 ;
        RECT 96.160 177.420 96.420 177.740 ;
        RECT 96.680 177.595 96.820 177.760 ;
        RECT 96.610 177.225 96.890 177.595 ;
        RECT 96.620 176.740 96.880 177.060 ;
        RECT 96.680 175.360 96.820 176.740 ;
        RECT 98.980 175.440 99.120 182.180 ;
        RECT 100.360 181.820 100.500 183.200 ;
        RECT 100.300 181.500 100.560 181.820 ;
        RECT 100.820 180.800 100.960 184.560 ;
        RECT 101.680 182.180 101.940 182.500 ;
        RECT 101.740 180.800 101.880 182.180 ;
        RECT 102.200 182.160 102.340 185.240 ;
        RECT 103.060 184.220 103.320 184.540 ;
        RECT 103.980 184.220 104.240 184.540 ;
        RECT 102.600 182.520 102.860 182.840 ;
        RECT 102.140 181.840 102.400 182.160 ;
        RECT 100.760 180.480 101.020 180.800 ;
        RECT 101.680 180.480 101.940 180.800 ;
        RECT 102.200 180.120 102.340 181.840 ;
        RECT 102.140 179.800 102.400 180.120 ;
        RECT 99.840 179.460 100.100 179.780 ;
        RECT 102.660 179.520 102.800 182.520 ;
        RECT 99.380 177.420 99.640 177.740 ;
        RECT 99.440 176.380 99.580 177.420 ;
        RECT 99.900 177.060 100.040 179.460 ;
        RECT 102.200 179.380 102.800 179.520 ;
        RECT 100.300 178.780 100.560 179.100 ;
        RECT 100.760 178.780 101.020 179.100 ;
        RECT 100.360 177.060 100.500 178.780 ;
        RECT 99.840 176.740 100.100 177.060 ;
        RECT 100.300 176.740 100.560 177.060 ;
        RECT 99.380 176.060 99.640 176.380 ;
        RECT 96.620 175.040 96.880 175.360 ;
        RECT 98.980 175.300 100.500 175.440 ;
        RECT 99.840 174.360 100.100 174.680 ;
        RECT 98.460 173.680 98.720 174.000 ;
        RECT 98.000 172.320 98.260 172.640 ;
        RECT 98.060 169.240 98.200 172.320 ;
        RECT 98.520 171.960 98.660 173.680 ;
        RECT 99.900 173.660 100.040 174.360 ;
        RECT 100.360 173.660 100.500 175.300 ;
        RECT 99.840 173.340 100.100 173.660 ;
        RECT 100.300 173.340 100.560 173.660 ;
        RECT 98.460 171.640 98.720 171.960 ;
        RECT 98.920 171.640 99.180 171.960 ;
        RECT 98.980 169.920 99.120 171.640 ;
        RECT 99.900 171.280 100.040 173.340 ;
        RECT 99.840 170.960 100.100 171.280 ;
        RECT 100.300 170.960 100.560 171.280 ;
        RECT 98.920 169.600 99.180 169.920 ;
        RECT 100.360 169.240 100.500 170.960 ;
        RECT 95.700 168.920 95.960 169.240 ;
        RECT 98.000 168.920 98.260 169.240 ;
        RECT 100.300 168.920 100.560 169.240 ;
        RECT 95.240 163.140 95.500 163.460 ;
        RECT 92.020 160.420 92.280 160.740 ;
        RECT 95.760 160.480 95.900 168.920 ;
        RECT 100.300 167.900 100.560 168.220 ;
        RECT 96.160 166.200 96.420 166.520 ;
        RECT 96.220 162.780 96.360 166.200 ;
        RECT 99.370 165.665 99.650 166.035 ;
        RECT 96.620 165.180 96.880 165.500 ;
        RECT 96.680 164.480 96.820 165.180 ;
        RECT 96.620 164.160 96.880 164.480 ;
        RECT 99.440 162.780 99.580 165.665 ;
        RECT 96.160 162.460 96.420 162.780 ;
        RECT 98.460 162.460 98.720 162.780 ;
        RECT 99.380 162.460 99.640 162.780 ;
        RECT 98.520 161.760 98.660 162.460 ;
        RECT 98.460 161.440 98.720 161.760 ;
        RECT 100.360 161.420 100.500 167.900 ;
        RECT 100.300 161.100 100.560 161.420 ;
        RECT 96.160 160.480 96.420 160.740 ;
        RECT 95.760 160.420 96.420 160.480 ;
        RECT 95.760 160.340 96.360 160.420 ;
        RECT 95.760 159.040 95.900 160.340 ;
        RECT 100.820 159.040 100.960 178.780 ;
        RECT 102.200 177.400 102.340 179.380 ;
        RECT 102.600 178.780 102.860 179.100 ;
        RECT 102.140 177.080 102.400 177.400 ;
        RECT 102.660 174.680 102.800 178.780 ;
        RECT 103.120 176.380 103.260 184.220 ;
        RECT 103.520 181.840 103.780 182.160 ;
        RECT 103.580 177.400 103.720 181.840 ;
        RECT 103.520 177.080 103.780 177.400 ;
        RECT 103.060 176.060 103.320 176.380 ;
        RECT 101.680 174.360 101.940 174.680 ;
        RECT 102.600 174.360 102.860 174.680 ;
        RECT 103.060 174.360 103.320 174.680 ;
        RECT 101.740 172.300 101.880 174.360 ;
        RECT 101.680 171.980 101.940 172.300 ;
        RECT 103.120 170.680 103.260 174.360 ;
        RECT 104.040 172.640 104.180 184.220 ;
        RECT 106.800 182.840 106.940 185.240 ;
        RECT 109.960 184.560 110.220 184.880 ;
        RECT 108.120 184.220 108.380 184.540 ;
        RECT 109.500 184.220 109.760 184.540 ;
        RECT 108.180 183.180 108.320 184.220 ;
        RECT 108.120 182.860 108.380 183.180 ;
        RECT 106.740 182.520 107.000 182.840 ;
        RECT 108.580 182.520 108.840 182.840 ;
        RECT 107.660 181.500 107.920 181.820 ;
        RECT 107.720 179.780 107.860 181.500 ;
        RECT 108.640 179.780 108.780 182.520 ;
        RECT 109.040 182.180 109.300 182.500 ;
        RECT 107.660 179.460 107.920 179.780 ;
        RECT 108.580 179.460 108.840 179.780 ;
        RECT 104.440 178.780 104.700 179.100 ;
        RECT 108.580 178.780 108.840 179.100 ;
        RECT 104.500 177.060 104.640 178.780 ;
        RECT 104.900 177.080 105.160 177.400 ;
        RECT 104.440 176.740 104.700 177.060 ;
        RECT 104.440 176.060 104.700 176.380 ;
        RECT 104.500 174.680 104.640 176.060 ;
        RECT 104.440 174.360 104.700 174.680 ;
        RECT 103.980 172.320 104.240 172.640 ;
        RECT 103.120 170.540 103.720 170.680 ;
        RECT 103.580 169.920 103.720 170.540 ;
        RECT 103.520 169.600 103.780 169.920 ;
        RECT 101.220 168.920 101.480 169.240 ;
        RECT 101.280 163.800 101.420 168.920 ;
        RECT 101.680 168.580 101.940 168.900 ;
        RECT 102.600 168.580 102.860 168.900 ;
        RECT 101.740 166.520 101.880 168.580 ;
        RECT 102.660 168.220 102.800 168.580 ;
        RECT 102.600 167.900 102.860 168.220 ;
        RECT 102.660 167.200 102.800 167.900 ;
        RECT 104.040 167.200 104.180 172.320 ;
        RECT 104.500 172.300 104.640 174.360 ;
        RECT 104.960 173.660 105.100 177.080 ;
        RECT 108.640 176.915 108.780 178.780 ;
        RECT 108.570 176.545 108.850 176.915 ;
        RECT 109.100 174.340 109.240 182.180 ;
        RECT 109.560 180.120 109.700 184.220 ;
        RECT 109.500 179.800 109.760 180.120 ;
        RECT 110.020 178.080 110.160 184.560 ;
        RECT 109.960 177.760 110.220 178.080 ;
        RECT 110.480 177.480 110.620 185.580 ;
        RECT 112.260 185.240 112.520 185.560 ;
        RECT 110.020 177.340 110.620 177.480 ;
        RECT 112.320 177.400 112.460 185.240 ;
        RECT 113.180 184.220 113.440 184.540 ;
        RECT 113.240 183.520 113.380 184.220 ;
        RECT 113.180 183.200 113.440 183.520 ;
        RECT 109.500 174.360 109.760 174.680 ;
        RECT 108.580 174.020 108.840 174.340 ;
        RECT 109.040 174.020 109.300 174.340 ;
        RECT 105.820 173.680 106.080 174.000 ;
        RECT 104.900 173.340 105.160 173.660 ;
        RECT 104.440 171.980 104.700 172.300 ;
        RECT 104.890 171.785 105.170 172.155 ;
        RECT 104.900 171.640 105.160 171.785 ;
        RECT 104.960 171.360 105.100 171.640 ;
        RECT 104.500 171.220 105.100 171.360 ;
        RECT 102.600 166.880 102.860 167.200 ;
        RECT 103.980 166.880 104.240 167.200 ;
        RECT 102.660 166.600 102.800 166.880 ;
        RECT 104.500 166.600 104.640 171.220 ;
        RECT 105.880 170.940 106.020 173.680 ;
        RECT 108.640 172.640 108.780 174.020 ;
        RECT 109.560 172.835 109.700 174.360 ;
        RECT 108.580 172.320 108.840 172.640 ;
        RECT 109.490 172.465 109.770 172.835 ;
        RECT 109.500 171.870 109.760 171.960 ;
        RECT 110.020 171.870 110.160 177.340 ;
        RECT 112.260 177.080 112.520 177.400 ;
        RECT 111.340 176.740 111.600 177.060 ;
        RECT 109.100 171.730 110.160 171.870 ;
        RECT 104.900 170.620 105.160 170.940 ;
        RECT 105.820 170.620 106.080 170.940 ;
        RECT 104.960 169.580 105.100 170.620 ;
        RECT 104.900 169.260 105.160 169.580 ;
        RECT 108.120 167.900 108.380 168.220 ;
        RECT 101.680 166.200 101.940 166.520 ;
        RECT 102.660 166.460 103.720 166.600 ;
        RECT 104.040 166.520 104.640 166.600 ;
        RECT 103.580 165.840 103.720 166.460 ;
        RECT 103.980 166.460 104.640 166.520 ;
        RECT 103.980 166.200 104.240 166.460 ;
        RECT 105.360 166.200 105.620 166.520 ;
        RECT 104.440 165.860 104.700 166.180 ;
        RECT 103.520 165.520 103.780 165.840 ;
        RECT 103.060 164.160 103.320 164.480 ;
        RECT 101.220 163.480 101.480 163.800 ;
        RECT 101.220 162.800 101.480 163.120 ;
        RECT 102.600 162.800 102.860 163.120 ;
        RECT 101.280 159.040 101.420 162.800 ;
        RECT 102.660 161.760 102.800 162.800 ;
        RECT 103.120 161.760 103.260 164.160 ;
        RECT 104.500 164.140 104.640 165.860 ;
        RECT 104.440 163.820 104.700 164.140 ;
        RECT 103.980 162.800 104.240 163.120 ;
        RECT 102.600 161.440 102.860 161.760 ;
        RECT 103.060 161.440 103.320 161.760 ;
        RECT 104.040 161.420 104.180 162.800 ;
        RECT 103.980 161.100 104.240 161.420 ;
        RECT 104.500 160.740 104.640 163.820 ;
        RECT 105.420 161.760 105.560 166.200 ;
        RECT 108.180 166.180 108.320 167.900 ;
        RECT 108.120 165.860 108.380 166.180 ;
        RECT 105.820 163.995 106.080 164.140 ;
        RECT 105.810 163.625 106.090 163.995 ;
        RECT 107.200 163.820 107.460 164.140 ;
        RECT 105.360 161.440 105.620 161.760 ;
        RECT 107.260 161.160 107.400 163.820 ;
        RECT 107.260 161.020 107.860 161.160 ;
        RECT 104.440 160.420 104.700 160.740 ;
        RECT 104.900 160.595 105.160 160.740 ;
        RECT 104.890 160.225 105.170 160.595 ;
        RECT 95.700 158.720 95.960 159.040 ;
        RECT 100.760 158.720 101.020 159.040 ;
        RECT 101.220 158.720 101.480 159.040 ;
        RECT 107.720 158.020 107.860 161.020 ;
        RECT 108.180 159.040 108.320 165.860 ;
        RECT 109.100 162.780 109.240 171.730 ;
        RECT 109.500 171.640 109.760 171.730 ;
        RECT 109.490 171.105 109.770 171.475 ;
        RECT 109.560 169.240 109.700 171.105 ;
        RECT 109.960 170.620 110.220 170.940 ;
        RECT 109.500 168.920 109.760 169.240 ;
        RECT 109.560 167.200 109.700 168.920 ;
        RECT 110.020 168.220 110.160 170.620 ;
        RECT 109.960 167.900 110.220 168.220 ;
        RECT 109.500 166.880 109.760 167.200 ;
        RECT 110.880 166.200 111.140 166.520 ;
        RECT 109.960 165.180 110.220 165.500 ;
        RECT 110.020 163.460 110.160 165.180 ;
        RECT 109.960 163.140 110.220 163.460 ;
        RECT 109.040 162.460 109.300 162.780 ;
        RECT 110.940 161.760 111.080 166.200 ;
        RECT 111.400 165.840 111.540 176.740 ;
        RECT 112.320 174.680 112.460 177.080 ;
        RECT 112.260 174.360 112.520 174.680 ;
        RECT 113.240 173.660 113.380 183.200 ;
        RECT 113.640 179.800 113.900 180.120 ;
        RECT 111.800 173.340 112.060 173.660 ;
        RECT 113.180 173.340 113.440 173.660 ;
        RECT 111.860 167.960 112.000 173.340 ;
        RECT 112.260 169.435 112.520 169.580 ;
        RECT 112.250 169.065 112.530 169.435 ;
        RECT 111.860 167.820 112.460 167.960 ;
        RECT 111.800 166.540 112.060 166.860 ;
        RECT 111.340 165.520 111.600 165.840 ;
        RECT 110.880 161.440 111.140 161.760 ;
        RECT 108.580 160.080 108.840 160.400 ;
        RECT 108.120 158.720 108.380 159.040 ;
        RECT 108.640 158.700 108.780 160.080 ;
        RECT 111.860 159.040 112.000 166.540 ;
        RECT 112.320 161.760 112.460 167.820 ;
        RECT 112.260 161.440 112.520 161.760 ;
        RECT 111.800 158.720 112.060 159.040 ;
        RECT 108.580 158.380 108.840 158.700 ;
        RECT 43.720 157.930 43.980 158.020 ;
        RECT 48.780 157.930 49.040 158.020 ;
        RECT 43.320 157.790 43.980 157.930 ;
        RECT 43.320 155.950 43.460 157.790 ;
        RECT 43.720 157.700 43.980 157.790 ;
        RECT 48.380 157.790 49.040 157.930 ;
        RECT 48.380 155.950 48.520 157.790 ;
        RECT 48.780 157.700 49.040 157.790 ;
        RECT 53.380 157.700 53.640 158.020 ;
        RECT 58.900 157.700 59.160 158.020 ;
        RECT 63.960 157.700 64.220 158.020 ;
        RECT 69.940 157.700 70.200 158.020 ;
        RECT 74.080 157.700 74.340 158.020 ;
        RECT 75.920 157.700 76.180 158.020 ;
        RECT 76.380 157.700 76.640 158.020 ;
        RECT 80.060 157.700 80.320 158.020 ;
        RECT 89.260 157.700 89.520 158.020 ;
        RECT 91.560 157.700 91.820 158.020 ;
        RECT 94.320 157.700 94.580 158.020 ;
        RECT 99.380 157.700 99.640 158.020 ;
        RECT 104.440 157.700 104.700 158.020 ;
        RECT 107.660 157.700 107.920 158.020 ;
        RECT 109.040 157.700 109.300 158.020 ;
        RECT 53.440 155.950 53.580 157.700 ;
        RECT 58.960 156.400 59.100 157.700 ;
        RECT 64.020 156.400 64.160 157.700 ;
        RECT 58.500 156.260 59.100 156.400 ;
        RECT 63.560 156.260 64.160 156.400 ;
        RECT 68.620 156.260 69.220 156.400 ;
        RECT 58.500 155.950 58.640 156.260 ;
        RECT 63.560 155.950 63.700 156.260 ;
        RECT 68.620 155.950 68.760 156.260 ;
        RECT 43.250 136.540 43.530 155.950 ;
        RECT 36.810 136.260 43.530 136.540 ;
        RECT 36.810 130.880 37.095 136.260 ;
        RECT 48.310 135.540 48.590 155.950 ;
        RECT 38.410 135.260 48.590 135.540 ;
        RECT 38.410 130.890 38.690 135.260 ;
        RECT 53.370 134.540 53.650 155.950 ;
        RECT 58.430 136.540 58.710 155.950 ;
        RECT 63.490 136.540 63.770 155.950 ;
        RECT 58.430 136.260 59.190 136.540 ;
        RECT 40.010 134.260 53.650 134.540 ;
        RECT 40.010 130.890 40.295 134.260 ;
        RECT 38.060 130.885 39.060 130.890 ;
        RECT 36.465 129.880 37.470 130.880 ;
        RECT 38.060 129.890 39.065 130.885 ;
        RECT 39.670 130.880 40.670 130.890 ;
        RECT 58.905 130.880 59.190 136.260 ;
        RECT 60.460 136.260 63.770 136.540 ;
        RECT 60.460 130.885 60.750 136.260 ;
        RECT 68.550 135.540 68.830 155.950 ;
        RECT 69.080 155.720 69.220 156.260 ;
        RECT 70.000 155.720 70.140 157.700 ;
        RECT 74.140 156.400 74.280 157.700 ;
        RECT 73.680 156.260 74.280 156.400 ;
        RECT 80.120 156.320 80.260 157.700 ;
        RECT 83.740 157.360 84.000 157.680 ;
        RECT 73.680 155.950 73.820 156.260 ;
        RECT 79.140 156.230 79.400 156.320 ;
        RECT 78.740 156.090 79.400 156.230 ;
        RECT 78.740 155.950 78.880 156.090 ;
        RECT 79.140 156.000 79.400 156.090 ;
        RECT 80.060 156.000 80.320 156.320 ;
        RECT 83.800 155.950 83.940 157.360 ;
        RECT 89.320 156.400 89.460 157.700 ;
        RECT 94.380 156.400 94.520 157.700 ;
        RECT 99.440 156.400 99.580 157.700 ;
        RECT 104.500 156.400 104.640 157.700 ;
        RECT 88.860 156.260 89.460 156.400 ;
        RECT 93.920 156.260 94.520 156.400 ;
        RECT 98.980 156.260 99.580 156.400 ;
        RECT 104.040 156.260 104.640 156.400 ;
        RECT 88.860 155.950 89.000 156.260 ;
        RECT 93.920 155.950 94.060 156.260 ;
        RECT 98.980 155.950 99.120 156.260 ;
        RECT 104.040 155.950 104.180 156.260 ;
        RECT 109.100 155.950 109.240 157.700 ;
        RECT 113.700 157.680 113.840 179.800 ;
        RECT 114.560 173.340 114.820 173.660 ;
        RECT 114.100 157.700 114.360 158.020 ;
        RECT 113.640 157.360 113.900 157.680 ;
        RECT 114.160 155.950 114.300 157.700 ;
        RECT 114.620 157.340 114.760 173.340 ;
        RECT 117.380 167.820 117.520 187.280 ;
        RECT 116.920 167.680 117.520 167.820 ;
        RECT 116.920 164.480 117.060 167.680 ;
        RECT 116.860 164.160 117.120 164.480 ;
        RECT 114.560 157.020 114.820 157.340 ;
        RECT 69.080 155.580 70.140 155.720 ;
        RECT 62.110 135.425 68.830 135.540 ;
        RECT 62.100 135.260 68.830 135.425 ;
        RECT 60.125 130.880 61.125 130.885 ;
        RECT 62.100 130.880 62.390 135.260 ;
        RECT 73.610 134.540 73.890 155.950 ;
        RECT 78.670 136.540 78.950 155.950 ;
        RECT 83.730 136.540 84.010 155.950 ;
        RECT 78.670 136.260 81.840 136.540 ;
        RECT 63.660 134.260 73.890 134.540 ;
        RECT 63.660 130.890 63.945 134.260 ;
        RECT 63.320 130.885 64.320 130.890 ;
        RECT 38.065 129.885 39.065 129.890 ;
        RECT 39.665 129.890 40.670 130.880 ;
        RECT 36.840 106.880 37.090 129.880 ;
        RECT 38.440 129.510 38.690 129.885 ;
        RECT 39.665 129.880 40.665 129.890 ;
        RECT 58.525 129.880 59.530 130.880 ;
        RECT 60.125 129.885 61.130 130.880 ;
        RECT 60.130 129.880 61.130 129.885 ;
        RECT 61.720 129.880 62.725 130.880 ;
        RECT 63.320 129.890 64.325 130.885 ;
        RECT 81.560 130.880 81.840 136.260 ;
        RECT 83.160 136.260 84.010 136.540 ;
        RECT 83.160 130.885 83.440 136.260 ;
        RECT 88.790 135.540 89.070 155.950 ;
        RECT 84.760 135.260 89.070 135.540 ;
        RECT 82.785 130.880 83.785 130.885 ;
        RECT 84.760 130.880 85.040 135.260 ;
        RECT 93.850 134.540 94.130 155.950 ;
        RECT 86.360 134.260 94.130 134.540 ;
        RECT 98.910 134.540 99.190 155.950 ;
        RECT 103.970 135.540 104.250 155.950 ;
        RECT 109.030 135.540 109.310 155.950 ;
        RECT 103.970 135.260 106.090 135.540 ;
        RECT 98.910 134.260 104.490 134.540 ;
        RECT 86.360 130.885 86.640 134.260 ;
        RECT 85.985 130.880 86.985 130.885 ;
        RECT 104.210 130.880 104.490 134.260 ;
        RECT 105.810 130.885 106.090 135.260 ;
        RECT 107.410 135.260 109.310 135.540 ;
        RECT 105.445 130.880 106.445 130.885 ;
        RECT 107.410 130.880 107.690 135.260 ;
        RECT 114.090 134.540 114.370 155.950 ;
        RECT 109.010 134.260 114.370 134.540 ;
        RECT 109.010 130.885 109.290 134.260 ;
        RECT 108.645 130.880 109.645 130.885 ;
        RECT 63.325 129.885 64.325 129.890 ;
        RECT 37.450 129.260 38.690 129.510 ;
        RECT 37.450 128.920 37.695 129.260 ;
        RECT 40.040 129.010 40.290 129.880 ;
        RECT 37.445 128.445 37.695 128.920 ;
        RECT 37.440 128.070 37.695 128.445 ;
        RECT 38.040 128.760 40.290 129.010 ;
        RECT 36.800 105.820 37.130 106.880 ;
        RECT 34.840 102.940 35.840 103.940 ;
        RECT 37.440 89.540 37.690 128.070 ;
        RECT 37.400 88.480 37.730 89.540 ;
        RECT 34.840 85.600 35.840 86.600 ;
        RECT 38.040 72.200 38.290 128.760 ;
        RECT 57.500 120.280 58.500 121.280 ;
        RECT 47.740 110.635 48.740 110.670 ;
        RECT 49.620 110.635 50.620 110.670 ;
        RECT 51.500 110.635 52.500 110.670 ;
        RECT 40.230 110.590 41.220 110.630 ;
        RECT 42.100 110.590 43.080 110.630 ;
        RECT 40.230 110.340 43.080 110.590 ;
        RECT 47.740 110.385 52.500 110.635 ;
        RECT 47.740 110.350 48.740 110.385 ;
        RECT 49.620 110.350 50.620 110.385 ;
        RECT 51.500 110.350 52.500 110.385 ;
        RECT 40.230 110.310 41.220 110.340 ;
        RECT 42.100 110.310 43.080 110.340 ;
        RECT 53.230 109.285 54.230 109.400 ;
        RECT 43.565 109.035 54.230 109.285 ;
        RECT 40.240 107.770 41.200 108.030 ;
        RECT 42.120 107.770 43.090 108.030 ;
        RECT 40.240 107.520 43.090 107.770 ;
        RECT 40.240 107.260 41.200 107.520 ;
        RECT 42.120 107.250 43.090 107.520 ;
        RECT 43.565 106.865 43.815 109.035 ;
        RECT 44.360 108.600 53.030 108.840 ;
        RECT 44.360 108.030 44.600 108.600 ;
        RECT 45.145 108.180 47.420 108.420 ;
        RECT 44.000 107.260 44.960 108.030 ;
        RECT 43.565 106.615 44.050 106.865 ;
        RECT 43.800 105.710 44.050 106.615 ;
        RECT 39.820 105.100 40.420 105.710 ;
        RECT 43.620 105.110 44.230 105.710 ;
        RECT 39.990 104.675 40.240 105.100 ;
        RECT 43.800 104.675 44.050 105.110 ;
        RECT 39.990 104.425 44.050 104.675 ;
        RECT 39.990 103.940 40.240 104.425 ;
        RECT 43.800 103.940 44.050 104.425 ;
        RECT 38.590 102.940 40.590 103.940 ;
        RECT 43.620 103.340 44.230 103.940 ;
        RECT 44.370 102.690 44.610 107.260 ;
        RECT 45.145 106.860 45.705 108.180 ;
        RECT 45.880 107.260 46.840 108.030 ;
        RECT 40.600 102.450 44.610 102.690 ;
        RECT 46.250 104.680 46.490 107.260 ;
        RECT 47.180 105.520 47.420 108.180 ;
        RECT 47.740 107.770 48.740 108.030 ;
        RECT 49.620 107.770 50.620 108.030 ;
        RECT 51.500 107.770 52.500 108.030 ;
        RECT 47.740 107.520 52.500 107.770 ;
        RECT 52.790 107.880 53.030 108.600 ;
        RECT 53.230 108.400 54.230 109.035 ;
        RECT 53.230 107.880 54.230 108.100 ;
        RECT 52.790 107.640 54.230 107.880 ;
        RECT 47.740 107.260 48.740 107.520 ;
        RECT 49.620 107.260 50.620 107.520 ;
        RECT 51.500 107.260 52.500 107.520 ;
        RECT 53.230 107.100 54.230 107.640 ;
        RECT 53.230 106.445 54.230 106.820 ;
        RECT 54.570 106.445 54.820 110.670 ;
        RECT 55.040 107.440 55.300 107.760 ;
        RECT 53.230 106.330 54.820 106.445 ;
        RECT 49.430 106.195 54.820 106.330 ;
        RECT 49.430 106.090 54.230 106.195 ;
        RECT 48.590 105.520 49.190 105.710 ;
        RECT 47.180 105.280 49.190 105.520 ;
        RECT 48.590 105.110 49.190 105.280 ;
        RECT 49.430 104.680 49.670 106.090 ;
        RECT 53.230 105.820 54.230 106.090 ;
        RECT 50.470 105.110 51.070 105.710 ;
        RECT 46.250 104.440 49.670 104.680 ;
        RECT 40.600 99.740 40.840 102.450 ;
        RECT 46.250 101.640 46.490 104.440 ;
        RECT 50.645 104.010 50.895 105.110 ;
        RECT 48.580 103.830 49.190 104.010 ;
        RECT 42.480 101.400 46.490 101.640 ;
        RECT 47.220 103.590 49.190 103.830 ;
        RECT 40.240 98.980 41.200 99.740 ;
        RECT 41.410 98.540 41.940 100.180 ;
        RECT 42.480 99.740 42.720 101.400 ;
        RECT 42.130 98.980 43.070 99.740 ;
        RECT 44.000 99.485 44.960 99.750 ;
        RECT 45.880 99.485 46.840 99.750 ;
        RECT 44.000 99.235 46.840 99.485 ;
        RECT 44.000 98.970 44.960 99.235 ;
        RECT 45.880 98.970 46.840 99.235 ;
        RECT 41.555 98.260 41.795 98.540 ;
        RECT 47.220 98.260 47.460 103.590 ;
        RECT 48.580 103.410 49.190 103.590 ;
        RECT 50.460 103.410 51.070 104.010 ;
        RECT 47.740 99.485 48.740 99.750 ;
        RECT 49.620 99.485 50.620 99.750 ;
        RECT 47.740 99.235 50.620 99.485 ;
        RECT 47.740 98.970 48.740 99.235 ;
        RECT 49.620 98.970 50.620 99.235 ;
        RECT 41.555 98.020 47.460 98.260 ;
        RECT 44.000 94.240 46.840 94.560 ;
        RECT 47.740 93.295 48.740 93.330 ;
        RECT 49.620 93.295 50.620 93.330 ;
        RECT 51.500 93.295 52.500 93.330 ;
        RECT 40.230 93.250 41.220 93.290 ;
        RECT 42.100 93.250 43.080 93.290 ;
        RECT 40.230 93.000 43.080 93.250 ;
        RECT 47.740 93.045 52.500 93.295 ;
        RECT 47.740 93.010 48.740 93.045 ;
        RECT 49.620 93.010 50.620 93.045 ;
        RECT 51.500 93.010 52.500 93.045 ;
        RECT 40.230 92.970 41.220 93.000 ;
        RECT 42.100 92.970 43.080 93.000 ;
        RECT 53.230 91.945 54.230 92.060 ;
        RECT 43.565 91.695 54.230 91.945 ;
        RECT 40.240 90.430 41.200 90.690 ;
        RECT 42.120 90.430 43.090 90.690 ;
        RECT 40.240 90.180 43.090 90.430 ;
        RECT 40.240 89.920 41.200 90.180 ;
        RECT 42.120 89.910 43.090 90.180 ;
        RECT 43.565 89.525 43.815 91.695 ;
        RECT 44.360 91.260 53.030 91.500 ;
        RECT 44.360 90.690 44.600 91.260 ;
        RECT 45.145 90.840 47.420 91.080 ;
        RECT 44.000 89.920 44.960 90.690 ;
        RECT 43.565 89.275 44.050 89.525 ;
        RECT 43.800 88.370 44.050 89.275 ;
        RECT 39.820 87.760 40.420 88.370 ;
        RECT 43.620 87.770 44.230 88.370 ;
        RECT 39.990 87.335 40.240 87.760 ;
        RECT 43.800 87.335 44.050 87.770 ;
        RECT 39.990 87.085 44.050 87.335 ;
        RECT 39.990 86.600 40.240 87.085 ;
        RECT 43.800 86.600 44.050 87.085 ;
        RECT 38.590 85.600 40.590 86.600 ;
        RECT 43.620 86.000 44.230 86.600 ;
        RECT 44.370 85.350 44.610 89.920 ;
        RECT 45.145 89.520 45.705 90.840 ;
        RECT 45.880 89.920 46.840 90.690 ;
        RECT 40.600 85.110 44.610 85.350 ;
        RECT 46.250 87.340 46.490 89.920 ;
        RECT 47.180 88.180 47.420 90.840 ;
        RECT 47.740 90.430 48.740 90.690 ;
        RECT 49.620 90.430 50.620 90.690 ;
        RECT 51.500 90.430 52.500 90.690 ;
        RECT 47.740 90.180 52.500 90.430 ;
        RECT 52.790 90.540 53.030 91.260 ;
        RECT 53.230 91.060 54.230 91.695 ;
        RECT 53.230 90.540 54.230 90.760 ;
        RECT 52.790 90.300 54.230 90.540 ;
        RECT 47.740 89.920 48.740 90.180 ;
        RECT 49.620 89.920 50.620 90.180 ;
        RECT 51.500 89.920 52.500 90.180 ;
        RECT 53.230 89.760 54.230 90.300 ;
        RECT 53.230 89.105 54.230 89.480 ;
        RECT 54.570 89.105 54.820 106.195 ;
        RECT 55.045 102.335 55.295 107.440 ;
        RECT 56.220 102.750 56.570 104.970 ;
        RECT 57.500 102.940 58.500 103.940 ;
        RECT 56.270 102.335 56.520 102.750 ;
        RECT 55.045 102.085 56.520 102.335 ;
        RECT 56.270 101.680 56.520 102.085 ;
        RECT 56.220 99.460 56.570 101.680 ;
        RECT 56.220 94.960 56.570 97.180 ;
        RECT 56.270 92.130 56.520 94.960 ;
        RECT 55.040 90.100 55.300 90.420 ;
        RECT 53.230 88.990 54.820 89.105 ;
        RECT 49.430 88.855 54.820 88.990 ;
        RECT 49.430 88.750 54.230 88.855 ;
        RECT 48.590 88.180 49.190 88.370 ;
        RECT 47.180 87.940 49.190 88.180 ;
        RECT 48.590 87.770 49.190 87.940 ;
        RECT 49.430 87.340 49.670 88.750 ;
        RECT 53.230 88.480 54.230 88.750 ;
        RECT 50.470 87.770 51.070 88.370 ;
        RECT 46.250 87.100 49.670 87.340 ;
        RECT 40.600 82.400 40.840 85.110 ;
        RECT 46.250 84.300 46.490 87.100 ;
        RECT 50.645 86.670 50.895 87.770 ;
        RECT 48.580 86.490 49.190 86.670 ;
        RECT 42.480 84.060 46.490 84.300 ;
        RECT 47.220 86.250 49.190 86.490 ;
        RECT 40.240 81.640 41.200 82.400 ;
        RECT 41.410 81.200 41.940 82.840 ;
        RECT 42.480 82.400 42.720 84.060 ;
        RECT 42.130 81.640 43.070 82.400 ;
        RECT 44.000 82.145 44.960 82.410 ;
        RECT 45.880 82.145 46.840 82.410 ;
        RECT 44.000 81.895 46.840 82.145 ;
        RECT 44.000 81.630 44.960 81.895 ;
        RECT 45.880 81.630 46.840 81.895 ;
        RECT 41.555 80.920 41.795 81.200 ;
        RECT 47.220 80.920 47.460 86.250 ;
        RECT 48.580 86.070 49.190 86.250 ;
        RECT 50.460 86.070 51.070 86.670 ;
        RECT 47.740 82.145 48.740 82.410 ;
        RECT 49.620 82.145 50.620 82.410 ;
        RECT 47.740 81.895 50.620 82.145 ;
        RECT 47.740 81.630 48.740 81.895 ;
        RECT 49.620 81.630 50.620 81.895 ;
        RECT 41.555 80.680 47.460 80.920 ;
        RECT 44.000 76.900 46.840 77.220 ;
        RECT 47.740 75.955 48.740 75.990 ;
        RECT 49.620 75.955 50.620 75.990 ;
        RECT 51.500 75.955 52.500 75.990 ;
        RECT 40.230 75.910 41.220 75.950 ;
        RECT 42.100 75.910 43.080 75.950 ;
        RECT 40.230 75.660 43.080 75.910 ;
        RECT 47.740 75.705 52.500 75.955 ;
        RECT 47.740 75.670 48.740 75.705 ;
        RECT 49.620 75.670 50.620 75.705 ;
        RECT 51.500 75.670 52.500 75.705 ;
        RECT 40.230 75.630 41.220 75.660 ;
        RECT 42.100 75.630 43.080 75.660 ;
        RECT 53.230 74.605 54.230 74.720 ;
        RECT 43.565 74.355 54.230 74.605 ;
        RECT 40.240 73.090 41.200 73.350 ;
        RECT 42.120 73.090 43.090 73.350 ;
        RECT 40.240 72.840 43.090 73.090 ;
        RECT 40.240 72.580 41.200 72.840 ;
        RECT 42.120 72.570 43.090 72.840 ;
        RECT 38.000 71.140 38.330 72.200 ;
        RECT 43.565 72.185 43.815 74.355 ;
        RECT 44.360 73.920 53.030 74.160 ;
        RECT 44.360 73.350 44.600 73.920 ;
        RECT 45.145 73.500 47.420 73.740 ;
        RECT 44.000 72.580 44.960 73.350 ;
        RECT 43.565 71.935 44.050 72.185 ;
        RECT 43.800 71.030 44.050 71.935 ;
        RECT 39.820 70.420 40.420 71.030 ;
        RECT 43.620 70.430 44.230 71.030 ;
        RECT 39.990 69.995 40.240 70.420 ;
        RECT 43.800 69.995 44.050 70.430 ;
        RECT 39.990 69.745 44.050 69.995 ;
        RECT 39.990 69.260 40.240 69.745 ;
        RECT 43.800 69.260 44.050 69.745 ;
        RECT 34.840 68.260 35.840 69.260 ;
        RECT 38.590 68.260 40.590 69.260 ;
        RECT 43.620 68.660 44.230 69.260 ;
        RECT 44.370 68.010 44.610 72.580 ;
        RECT 45.145 72.180 45.705 73.500 ;
        RECT 45.880 72.580 46.840 73.350 ;
        RECT 40.600 67.770 44.610 68.010 ;
        RECT 46.250 70.000 46.490 72.580 ;
        RECT 47.180 70.840 47.420 73.500 ;
        RECT 47.740 73.090 48.740 73.350 ;
        RECT 49.620 73.090 50.620 73.350 ;
        RECT 51.500 73.090 52.500 73.350 ;
        RECT 47.740 72.840 52.500 73.090 ;
        RECT 52.790 73.200 53.030 73.920 ;
        RECT 53.230 73.720 54.230 74.355 ;
        RECT 53.230 73.200 54.230 73.420 ;
        RECT 52.790 72.960 54.230 73.200 ;
        RECT 47.740 72.580 48.740 72.840 ;
        RECT 49.620 72.580 50.620 72.840 ;
        RECT 51.500 72.580 52.500 72.840 ;
        RECT 53.230 72.420 54.230 72.960 ;
        RECT 53.230 71.765 54.230 72.140 ;
        RECT 54.570 71.765 54.820 88.855 ;
        RECT 55.045 84.995 55.295 90.100 ;
        RECT 56.220 89.910 56.570 92.130 ;
        RECT 56.220 85.410 56.570 87.630 ;
        RECT 57.500 85.600 58.500 86.600 ;
        RECT 56.270 84.995 56.520 85.410 ;
        RECT 55.045 84.745 56.520 84.995 ;
        RECT 56.270 84.340 56.520 84.745 ;
        RECT 56.220 82.120 56.570 84.340 ;
        RECT 56.220 77.620 56.570 79.840 ;
        RECT 56.270 74.790 56.520 77.620 ;
        RECT 55.040 72.760 55.300 73.080 ;
        RECT 53.230 71.650 54.820 71.765 ;
        RECT 49.430 71.515 54.820 71.650 ;
        RECT 49.430 71.410 54.230 71.515 ;
        RECT 48.590 70.840 49.190 71.030 ;
        RECT 47.180 70.600 49.190 70.840 ;
        RECT 48.590 70.430 49.190 70.600 ;
        RECT 49.430 70.000 49.670 71.410 ;
        RECT 53.230 71.140 54.230 71.410 ;
        RECT 50.470 70.430 51.070 71.030 ;
        RECT 46.250 69.760 49.670 70.000 ;
        RECT 40.600 65.060 40.840 67.770 ;
        RECT 46.250 66.960 46.490 69.760 ;
        RECT 50.645 69.330 50.895 70.430 ;
        RECT 48.580 69.150 49.190 69.330 ;
        RECT 42.480 66.720 46.490 66.960 ;
        RECT 47.220 68.910 49.190 69.150 ;
        RECT 40.240 64.300 41.200 65.060 ;
        RECT 41.410 63.860 41.940 65.500 ;
        RECT 42.480 65.060 42.720 66.720 ;
        RECT 42.130 64.300 43.070 65.060 ;
        RECT 44.000 64.805 44.960 65.070 ;
        RECT 45.880 64.805 46.840 65.070 ;
        RECT 44.000 64.555 46.840 64.805 ;
        RECT 44.000 64.290 44.960 64.555 ;
        RECT 45.880 64.290 46.840 64.555 ;
        RECT 41.555 63.580 41.795 63.860 ;
        RECT 47.220 63.580 47.460 68.910 ;
        RECT 48.580 68.730 49.190 68.910 ;
        RECT 50.460 68.730 51.070 69.330 ;
        RECT 47.740 64.805 48.740 65.070 ;
        RECT 49.620 64.805 50.620 65.070 ;
        RECT 47.740 64.555 50.620 64.805 ;
        RECT 47.740 64.290 48.740 64.555 ;
        RECT 49.620 64.290 50.620 64.555 ;
        RECT 41.555 63.340 47.460 63.580 ;
        RECT 44.000 59.560 46.840 59.880 ;
        RECT 54.570 58.455 54.820 71.515 ;
        RECT 55.045 67.655 55.295 72.760 ;
        RECT 56.220 72.570 56.570 74.790 ;
        RECT 58.900 72.200 59.150 129.880 ;
        RECT 60.500 129.510 60.750 129.880 ;
        RECT 59.505 129.260 60.750 129.510 ;
        RECT 59.505 128.475 59.755 129.260 ;
        RECT 62.100 129.010 62.350 129.880 ;
        RECT 59.500 128.070 59.755 128.475 ;
        RECT 60.100 128.760 62.350 129.010 ;
        RECT 59.500 89.540 59.750 128.070 ;
        RECT 60.100 106.880 60.350 128.760 ;
        RECT 63.700 128.510 63.950 129.885 ;
        RECT 81.180 129.880 82.185 130.880 ;
        RECT 82.780 129.885 83.785 130.880 ;
        RECT 82.780 129.880 83.780 129.885 ;
        RECT 84.385 129.880 85.390 130.880 ;
        RECT 85.980 129.885 86.985 130.880 ;
        RECT 85.980 129.880 86.980 129.885 ;
        RECT 103.840 129.880 104.845 130.880 ;
        RECT 105.440 129.885 106.445 130.880 ;
        RECT 105.440 129.880 106.440 129.885 ;
        RECT 107.040 129.880 108.045 130.880 ;
        RECT 108.645 129.885 109.650 130.880 ;
        RECT 108.650 129.880 109.650 129.885 ;
        RECT 60.700 128.260 63.950 128.510 ;
        RECT 78.940 128.310 79.200 128.630 ;
        RECT 60.700 124.220 60.950 128.260 ;
        RECT 78.945 128.010 79.195 128.310 ;
        RECT 70.400 127.975 71.400 128.010 ;
        RECT 72.280 127.975 73.280 128.010 ;
        RECT 74.160 127.975 75.160 128.010 ;
        RECT 62.890 127.930 63.880 127.970 ;
        RECT 64.760 127.930 65.740 127.970 ;
        RECT 62.890 127.680 65.740 127.930 ;
        RECT 70.400 127.725 75.160 127.975 ;
        RECT 70.400 127.690 71.400 127.725 ;
        RECT 72.280 127.690 73.280 127.725 ;
        RECT 74.160 127.690 75.160 127.725 ;
        RECT 62.890 127.650 63.880 127.680 ;
        RECT 64.760 127.650 65.740 127.680 ;
        RECT 75.890 126.625 76.890 126.740 ;
        RECT 66.225 126.375 76.890 126.625 ;
        RECT 62.900 125.110 63.860 125.370 ;
        RECT 64.780 125.110 65.750 125.370 ;
        RECT 62.900 124.860 65.750 125.110 ;
        RECT 62.900 124.600 63.860 124.860 ;
        RECT 64.780 124.590 65.750 124.860 ;
        RECT 60.660 123.160 60.990 124.220 ;
        RECT 66.225 124.205 66.475 126.375 ;
        RECT 67.020 125.940 75.690 126.180 ;
        RECT 67.020 125.370 67.260 125.940 ;
        RECT 67.805 125.520 70.080 125.760 ;
        RECT 66.660 124.600 67.620 125.370 ;
        RECT 66.225 123.955 66.710 124.205 ;
        RECT 66.460 123.050 66.710 123.955 ;
        RECT 62.480 122.440 63.080 123.050 ;
        RECT 66.280 122.450 66.890 123.050 ;
        RECT 62.650 122.015 62.900 122.440 ;
        RECT 66.460 122.015 66.710 122.450 ;
        RECT 62.650 121.765 66.710 122.015 ;
        RECT 62.650 121.280 62.900 121.765 ;
        RECT 66.460 121.280 66.710 121.765 ;
        RECT 61.250 120.280 63.250 121.280 ;
        RECT 66.280 120.680 66.890 121.280 ;
        RECT 67.030 120.030 67.270 124.600 ;
        RECT 67.805 124.200 68.365 125.520 ;
        RECT 68.540 124.600 69.500 125.370 ;
        RECT 63.260 119.790 67.270 120.030 ;
        RECT 68.910 122.020 69.150 124.600 ;
        RECT 69.840 122.860 70.080 125.520 ;
        RECT 70.400 125.110 71.400 125.370 ;
        RECT 72.280 125.110 73.280 125.370 ;
        RECT 74.160 125.110 75.160 125.370 ;
        RECT 70.400 124.860 75.160 125.110 ;
        RECT 75.450 125.220 75.690 125.940 ;
        RECT 75.890 125.740 76.890 126.375 ;
        RECT 75.890 125.220 76.890 125.440 ;
        RECT 75.450 124.980 76.890 125.220 ;
        RECT 70.400 124.600 71.400 124.860 ;
        RECT 72.280 124.600 73.280 124.860 ;
        RECT 74.160 124.600 75.160 124.860 ;
        RECT 75.890 124.440 76.890 124.980 ;
        RECT 75.890 123.785 76.890 124.160 ;
        RECT 77.230 123.785 77.480 128.010 ;
        RECT 78.930 127.655 79.195 128.010 ;
        RECT 78.930 126.810 79.180 127.655 ;
        RECT 77.700 124.780 77.960 125.100 ;
        RECT 75.890 123.670 77.480 123.785 ;
        RECT 72.090 123.535 77.480 123.670 ;
        RECT 72.090 123.430 76.890 123.535 ;
        RECT 71.250 122.860 71.850 123.050 ;
        RECT 69.840 122.620 71.850 122.860 ;
        RECT 71.250 122.450 71.850 122.620 ;
        RECT 72.090 122.020 72.330 123.430 ;
        RECT 75.890 123.160 76.890 123.430 ;
        RECT 73.130 122.450 73.730 123.050 ;
        RECT 68.910 121.780 72.330 122.020 ;
        RECT 63.260 117.080 63.500 119.790 ;
        RECT 68.910 118.980 69.150 121.780 ;
        RECT 73.305 121.350 73.555 122.450 ;
        RECT 71.240 121.170 71.850 121.350 ;
        RECT 65.140 118.740 69.150 118.980 ;
        RECT 69.880 120.930 71.850 121.170 ;
        RECT 62.900 116.320 63.860 117.080 ;
        RECT 64.070 115.880 64.600 117.520 ;
        RECT 65.140 117.080 65.380 118.740 ;
        RECT 64.790 116.320 65.730 117.080 ;
        RECT 66.660 116.825 67.620 117.090 ;
        RECT 68.540 116.825 69.500 117.090 ;
        RECT 66.660 116.575 69.500 116.825 ;
        RECT 66.660 116.310 67.620 116.575 ;
        RECT 68.540 116.310 69.500 116.575 ;
        RECT 64.215 115.600 64.455 115.880 ;
        RECT 69.880 115.600 70.120 120.930 ;
        RECT 71.240 120.750 71.850 120.930 ;
        RECT 73.120 120.750 73.730 121.350 ;
        RECT 70.400 116.825 71.400 117.090 ;
        RECT 72.280 116.825 73.280 117.090 ;
        RECT 70.400 116.575 73.280 116.825 ;
        RECT 70.400 116.310 71.400 116.575 ;
        RECT 72.280 116.310 73.280 116.575 ;
        RECT 64.215 115.360 70.120 115.600 ;
        RECT 66.660 111.580 69.500 111.900 ;
        RECT 70.400 110.635 71.400 110.670 ;
        RECT 72.280 110.635 73.280 110.670 ;
        RECT 74.160 110.635 75.160 110.670 ;
        RECT 62.890 110.590 63.880 110.630 ;
        RECT 64.760 110.590 65.740 110.630 ;
        RECT 62.890 110.340 65.740 110.590 ;
        RECT 70.400 110.385 75.160 110.635 ;
        RECT 70.400 110.350 71.400 110.385 ;
        RECT 72.280 110.350 73.280 110.385 ;
        RECT 74.160 110.350 75.160 110.385 ;
        RECT 62.890 110.310 63.880 110.340 ;
        RECT 64.760 110.310 65.740 110.340 ;
        RECT 75.890 109.285 76.890 109.400 ;
        RECT 66.225 109.035 76.890 109.285 ;
        RECT 62.900 107.770 63.860 108.030 ;
        RECT 64.780 107.770 65.750 108.030 ;
        RECT 62.900 107.520 65.750 107.770 ;
        RECT 62.900 107.260 63.860 107.520 ;
        RECT 64.780 107.250 65.750 107.520 ;
        RECT 60.060 105.820 60.390 106.880 ;
        RECT 66.225 106.865 66.475 109.035 ;
        RECT 67.020 108.600 75.690 108.840 ;
        RECT 67.020 108.030 67.260 108.600 ;
        RECT 67.805 108.180 70.080 108.420 ;
        RECT 66.660 107.260 67.620 108.030 ;
        RECT 66.225 106.615 66.710 106.865 ;
        RECT 66.460 105.710 66.710 106.615 ;
        RECT 62.480 105.100 63.080 105.710 ;
        RECT 66.280 105.110 66.890 105.710 ;
        RECT 62.650 104.675 62.900 105.100 ;
        RECT 66.460 104.675 66.710 105.110 ;
        RECT 62.650 104.425 66.710 104.675 ;
        RECT 62.650 103.940 62.900 104.425 ;
        RECT 66.460 103.940 66.710 104.425 ;
        RECT 61.250 102.940 63.250 103.940 ;
        RECT 66.280 103.340 66.890 103.940 ;
        RECT 67.030 102.690 67.270 107.260 ;
        RECT 67.805 106.860 68.365 108.180 ;
        RECT 68.540 107.260 69.500 108.030 ;
        RECT 63.260 102.450 67.270 102.690 ;
        RECT 68.910 104.680 69.150 107.260 ;
        RECT 69.840 105.520 70.080 108.180 ;
        RECT 70.400 107.770 71.400 108.030 ;
        RECT 72.280 107.770 73.280 108.030 ;
        RECT 74.160 107.770 75.160 108.030 ;
        RECT 70.400 107.520 75.160 107.770 ;
        RECT 75.450 107.880 75.690 108.600 ;
        RECT 75.890 108.400 76.890 109.035 ;
        RECT 75.890 107.880 76.890 108.100 ;
        RECT 75.450 107.640 76.890 107.880 ;
        RECT 70.400 107.260 71.400 107.520 ;
        RECT 72.280 107.260 73.280 107.520 ;
        RECT 74.160 107.260 75.160 107.520 ;
        RECT 75.890 107.100 76.890 107.640 ;
        RECT 75.890 106.445 76.890 106.820 ;
        RECT 77.230 106.445 77.480 123.535 ;
        RECT 77.705 119.675 77.955 124.780 ;
        RECT 78.880 124.590 79.230 126.810 ;
        RECT 81.560 124.220 81.810 129.880 ;
        RECT 83.160 129.510 83.410 129.880 ;
        RECT 82.170 129.260 83.410 129.510 ;
        RECT 82.170 129.240 82.415 129.260 ;
        RECT 82.165 128.645 82.415 129.240 ;
        RECT 84.760 129.010 85.010 129.880 ;
        RECT 82.160 127.565 82.415 128.645 ;
        RECT 82.760 128.760 85.010 129.010 ;
        RECT 81.520 123.160 81.850 124.220 ;
        RECT 78.880 120.090 79.230 122.310 ;
        RECT 80.160 120.280 81.160 121.280 ;
        RECT 78.930 119.675 79.180 120.090 ;
        RECT 77.705 119.425 79.180 119.675 ;
        RECT 78.930 119.020 79.180 119.425 ;
        RECT 78.880 116.800 79.230 119.020 ;
        RECT 78.880 112.300 79.230 114.520 ;
        RECT 78.930 109.470 79.180 112.300 ;
        RECT 77.700 107.440 77.960 107.760 ;
        RECT 75.890 106.330 77.480 106.445 ;
        RECT 72.090 106.195 77.480 106.330 ;
        RECT 72.090 106.090 76.890 106.195 ;
        RECT 71.250 105.520 71.850 105.710 ;
        RECT 69.840 105.280 71.850 105.520 ;
        RECT 71.250 105.110 71.850 105.280 ;
        RECT 72.090 104.680 72.330 106.090 ;
        RECT 75.890 105.820 76.890 106.090 ;
        RECT 73.130 105.110 73.730 105.710 ;
        RECT 68.910 104.440 72.330 104.680 ;
        RECT 63.260 99.740 63.500 102.450 ;
        RECT 68.910 101.640 69.150 104.440 ;
        RECT 73.305 104.010 73.555 105.110 ;
        RECT 71.240 103.830 71.850 104.010 ;
        RECT 65.140 101.400 69.150 101.640 ;
        RECT 69.880 103.590 71.850 103.830 ;
        RECT 62.900 98.980 63.860 99.740 ;
        RECT 64.070 98.540 64.600 100.180 ;
        RECT 65.140 99.740 65.380 101.400 ;
        RECT 64.790 98.980 65.730 99.740 ;
        RECT 66.660 99.485 67.620 99.750 ;
        RECT 68.540 99.485 69.500 99.750 ;
        RECT 66.660 99.235 69.500 99.485 ;
        RECT 66.660 98.970 67.620 99.235 ;
        RECT 68.540 98.970 69.500 99.235 ;
        RECT 64.215 98.260 64.455 98.540 ;
        RECT 69.880 98.260 70.120 103.590 ;
        RECT 71.240 103.410 71.850 103.590 ;
        RECT 73.120 103.410 73.730 104.010 ;
        RECT 70.400 99.485 71.400 99.750 ;
        RECT 72.280 99.485 73.280 99.750 ;
        RECT 70.400 99.235 73.280 99.485 ;
        RECT 70.400 98.970 71.400 99.235 ;
        RECT 72.280 98.970 73.280 99.235 ;
        RECT 64.215 98.020 70.120 98.260 ;
        RECT 66.660 94.240 69.500 94.560 ;
        RECT 70.400 93.295 71.400 93.330 ;
        RECT 72.280 93.295 73.280 93.330 ;
        RECT 74.160 93.295 75.160 93.330 ;
        RECT 62.890 93.250 63.880 93.290 ;
        RECT 64.760 93.250 65.740 93.290 ;
        RECT 62.890 93.000 65.740 93.250 ;
        RECT 70.400 93.045 75.160 93.295 ;
        RECT 70.400 93.010 71.400 93.045 ;
        RECT 72.280 93.010 73.280 93.045 ;
        RECT 74.160 93.010 75.160 93.045 ;
        RECT 62.890 92.970 63.880 93.000 ;
        RECT 64.760 92.970 65.740 93.000 ;
        RECT 75.890 91.945 76.890 92.060 ;
        RECT 66.225 91.695 76.890 91.945 ;
        RECT 62.900 90.430 63.860 90.690 ;
        RECT 64.780 90.430 65.750 90.690 ;
        RECT 62.900 90.180 65.750 90.430 ;
        RECT 62.900 89.920 63.860 90.180 ;
        RECT 64.780 89.910 65.750 90.180 ;
        RECT 59.460 88.480 59.790 89.540 ;
        RECT 66.225 89.525 66.475 91.695 ;
        RECT 67.020 91.260 75.690 91.500 ;
        RECT 67.020 90.690 67.260 91.260 ;
        RECT 67.805 90.840 70.080 91.080 ;
        RECT 66.660 89.920 67.620 90.690 ;
        RECT 66.225 89.275 66.710 89.525 ;
        RECT 66.460 88.370 66.710 89.275 ;
        RECT 62.480 87.760 63.080 88.370 ;
        RECT 66.280 87.770 66.890 88.370 ;
        RECT 62.650 87.335 62.900 87.760 ;
        RECT 66.460 87.335 66.710 87.770 ;
        RECT 62.650 87.085 66.710 87.335 ;
        RECT 62.650 86.600 62.900 87.085 ;
        RECT 66.460 86.600 66.710 87.085 ;
        RECT 61.250 85.600 63.250 86.600 ;
        RECT 66.280 86.000 66.890 86.600 ;
        RECT 67.030 85.350 67.270 89.920 ;
        RECT 67.805 89.520 68.365 90.840 ;
        RECT 68.540 89.920 69.500 90.690 ;
        RECT 63.260 85.110 67.270 85.350 ;
        RECT 68.910 87.340 69.150 89.920 ;
        RECT 69.840 88.180 70.080 90.840 ;
        RECT 70.400 90.430 71.400 90.690 ;
        RECT 72.280 90.430 73.280 90.690 ;
        RECT 74.160 90.430 75.160 90.690 ;
        RECT 70.400 90.180 75.160 90.430 ;
        RECT 75.450 90.540 75.690 91.260 ;
        RECT 75.890 91.060 76.890 91.695 ;
        RECT 75.890 90.540 76.890 90.760 ;
        RECT 75.450 90.300 76.890 90.540 ;
        RECT 70.400 89.920 71.400 90.180 ;
        RECT 72.280 89.920 73.280 90.180 ;
        RECT 74.160 89.920 75.160 90.180 ;
        RECT 75.890 89.760 76.890 90.300 ;
        RECT 75.890 89.105 76.890 89.480 ;
        RECT 77.230 89.105 77.480 106.195 ;
        RECT 77.705 102.335 77.955 107.440 ;
        RECT 78.880 107.250 79.230 109.470 ;
        RECT 82.160 106.880 82.410 127.565 ;
        RECT 82.120 105.820 82.450 106.880 ;
        RECT 78.880 102.750 79.230 104.970 ;
        RECT 80.160 102.940 81.160 103.940 ;
        RECT 78.930 102.335 79.180 102.750 ;
        RECT 77.705 102.085 79.180 102.335 ;
        RECT 78.930 101.680 79.180 102.085 ;
        RECT 78.880 99.460 79.230 101.680 ;
        RECT 78.880 94.960 79.230 97.180 ;
        RECT 78.930 92.130 79.180 94.960 ;
        RECT 77.700 90.100 77.960 90.420 ;
        RECT 75.890 88.990 77.480 89.105 ;
        RECT 72.090 88.855 77.480 88.990 ;
        RECT 72.090 88.750 76.890 88.855 ;
        RECT 71.250 88.180 71.850 88.370 ;
        RECT 69.840 87.940 71.850 88.180 ;
        RECT 71.250 87.770 71.850 87.940 ;
        RECT 72.090 87.340 72.330 88.750 ;
        RECT 75.890 88.480 76.890 88.750 ;
        RECT 73.130 87.770 73.730 88.370 ;
        RECT 68.910 87.100 72.330 87.340 ;
        RECT 63.260 82.400 63.500 85.110 ;
        RECT 68.910 84.300 69.150 87.100 ;
        RECT 73.305 86.670 73.555 87.770 ;
        RECT 71.240 86.490 71.850 86.670 ;
        RECT 65.140 84.060 69.150 84.300 ;
        RECT 69.880 86.250 71.850 86.490 ;
        RECT 62.900 81.640 63.860 82.400 ;
        RECT 64.070 81.200 64.600 82.840 ;
        RECT 65.140 82.400 65.380 84.060 ;
        RECT 64.790 81.640 65.730 82.400 ;
        RECT 66.660 82.145 67.620 82.410 ;
        RECT 68.540 82.145 69.500 82.410 ;
        RECT 66.660 81.895 69.500 82.145 ;
        RECT 66.660 81.630 67.620 81.895 ;
        RECT 68.540 81.630 69.500 81.895 ;
        RECT 64.215 80.920 64.455 81.200 ;
        RECT 69.880 80.920 70.120 86.250 ;
        RECT 71.240 86.070 71.850 86.250 ;
        RECT 73.120 86.070 73.730 86.670 ;
        RECT 70.400 82.145 71.400 82.410 ;
        RECT 72.280 82.145 73.280 82.410 ;
        RECT 70.400 81.895 73.280 82.145 ;
        RECT 70.400 81.630 71.400 81.895 ;
        RECT 72.280 81.630 73.280 81.895 ;
        RECT 64.215 80.680 70.120 80.920 ;
        RECT 66.660 76.900 69.500 77.220 ;
        RECT 70.400 75.955 71.400 75.990 ;
        RECT 72.280 75.955 73.280 75.990 ;
        RECT 74.160 75.955 75.160 75.990 ;
        RECT 62.890 75.910 63.880 75.950 ;
        RECT 64.760 75.910 65.740 75.950 ;
        RECT 62.890 75.660 65.740 75.910 ;
        RECT 70.400 75.705 75.160 75.955 ;
        RECT 70.400 75.670 71.400 75.705 ;
        RECT 72.280 75.670 73.280 75.705 ;
        RECT 74.160 75.670 75.160 75.705 ;
        RECT 62.890 75.630 63.880 75.660 ;
        RECT 64.760 75.630 65.740 75.660 ;
        RECT 75.890 74.605 76.890 74.720 ;
        RECT 66.225 74.355 76.890 74.605 ;
        RECT 62.900 73.090 63.860 73.350 ;
        RECT 64.780 73.090 65.750 73.350 ;
        RECT 62.900 72.840 65.750 73.090 ;
        RECT 62.900 72.580 63.860 72.840 ;
        RECT 64.780 72.570 65.750 72.840 ;
        RECT 58.860 71.140 59.190 72.200 ;
        RECT 66.225 72.185 66.475 74.355 ;
        RECT 67.020 73.920 75.690 74.160 ;
        RECT 67.020 73.350 67.260 73.920 ;
        RECT 67.805 73.500 70.080 73.740 ;
        RECT 66.660 72.580 67.620 73.350 ;
        RECT 66.225 71.935 66.710 72.185 ;
        RECT 66.460 71.030 66.710 71.935 ;
        RECT 62.480 70.420 63.080 71.030 ;
        RECT 66.280 70.430 66.890 71.030 ;
        RECT 56.220 68.070 56.570 70.290 ;
        RECT 62.650 69.995 62.900 70.420 ;
        RECT 66.460 69.995 66.710 70.430 ;
        RECT 62.650 69.745 66.710 69.995 ;
        RECT 62.650 69.260 62.900 69.745 ;
        RECT 66.460 69.260 66.710 69.745 ;
        RECT 57.500 68.260 58.500 69.260 ;
        RECT 61.250 68.260 63.250 69.260 ;
        RECT 66.280 68.660 66.890 69.260 ;
        RECT 56.270 67.655 56.520 68.070 ;
        RECT 67.030 68.010 67.270 72.580 ;
        RECT 67.805 72.180 68.365 73.500 ;
        RECT 68.540 72.580 69.500 73.350 ;
        RECT 55.045 67.405 56.520 67.655 ;
        RECT 56.270 67.000 56.520 67.405 ;
        RECT 63.260 67.770 67.270 68.010 ;
        RECT 68.910 70.000 69.150 72.580 ;
        RECT 69.840 70.840 70.080 73.500 ;
        RECT 70.400 73.090 71.400 73.350 ;
        RECT 72.280 73.090 73.280 73.350 ;
        RECT 74.160 73.090 75.160 73.350 ;
        RECT 70.400 72.840 75.160 73.090 ;
        RECT 75.450 73.200 75.690 73.920 ;
        RECT 75.890 73.720 76.890 74.355 ;
        RECT 75.890 73.200 76.890 73.420 ;
        RECT 75.450 72.960 76.890 73.200 ;
        RECT 70.400 72.580 71.400 72.840 ;
        RECT 72.280 72.580 73.280 72.840 ;
        RECT 74.160 72.580 75.160 72.840 ;
        RECT 75.890 72.420 76.890 72.960 ;
        RECT 75.890 71.765 76.890 72.140 ;
        RECT 77.230 71.765 77.480 88.855 ;
        RECT 77.705 84.995 77.955 90.100 ;
        RECT 78.880 89.910 79.230 92.130 ;
        RECT 82.760 89.540 83.010 128.760 ;
        RECT 86.360 128.510 86.610 129.880 ;
        RECT 83.360 128.260 86.610 128.510 ;
        RECT 101.585 128.310 101.845 128.630 ;
        RECT 82.720 88.480 83.050 89.540 ;
        RECT 78.880 85.410 79.230 87.630 ;
        RECT 80.160 85.600 81.160 86.600 ;
        RECT 78.930 84.995 79.180 85.410 ;
        RECT 77.705 84.745 79.180 84.995 ;
        RECT 78.930 84.340 79.180 84.745 ;
        RECT 78.880 82.120 79.230 84.340 ;
        RECT 78.880 77.620 79.230 79.840 ;
        RECT 78.930 74.790 79.180 77.620 ;
        RECT 77.700 72.760 77.960 73.080 ;
        RECT 75.890 71.650 77.480 71.765 ;
        RECT 72.090 71.515 77.480 71.650 ;
        RECT 72.090 71.410 76.890 71.515 ;
        RECT 71.250 70.840 71.850 71.030 ;
        RECT 69.840 70.600 71.850 70.840 ;
        RECT 71.250 70.430 71.850 70.600 ;
        RECT 72.090 70.000 72.330 71.410 ;
        RECT 75.890 71.140 76.890 71.410 ;
        RECT 73.130 70.430 73.730 71.030 ;
        RECT 68.910 69.760 72.330 70.000 ;
        RECT 56.220 64.780 56.570 67.000 ;
        RECT 63.260 65.060 63.500 67.770 ;
        RECT 68.910 66.960 69.150 69.760 ;
        RECT 73.305 69.330 73.555 70.430 ;
        RECT 71.240 69.150 71.850 69.330 ;
        RECT 65.140 66.720 69.150 66.960 ;
        RECT 69.880 68.910 71.850 69.150 ;
        RECT 62.900 64.300 63.860 65.060 ;
        RECT 64.070 63.860 64.600 65.500 ;
        RECT 65.140 65.060 65.380 66.720 ;
        RECT 64.790 64.300 65.730 65.060 ;
        RECT 66.660 64.805 67.620 65.070 ;
        RECT 68.540 64.805 69.500 65.070 ;
        RECT 66.660 64.555 69.500 64.805 ;
        RECT 66.660 64.290 67.620 64.555 ;
        RECT 68.540 64.290 69.500 64.555 ;
        RECT 64.215 63.580 64.455 63.860 ;
        RECT 69.880 63.580 70.120 68.910 ;
        RECT 71.240 68.730 71.850 68.910 ;
        RECT 73.120 68.730 73.730 69.330 ;
        RECT 70.400 64.805 71.400 65.070 ;
        RECT 72.280 64.805 73.280 65.070 ;
        RECT 70.400 64.555 73.280 64.805 ;
        RECT 70.400 64.290 71.400 64.555 ;
        RECT 72.280 64.290 73.280 64.555 ;
        RECT 64.215 63.340 70.120 63.580 ;
        RECT 56.220 60.280 56.570 62.500 ;
        RECT 56.270 59.465 56.520 60.280 ;
        RECT 66.660 59.560 69.500 59.880 ;
        RECT 77.230 59.465 77.480 71.515 ;
        RECT 77.705 67.655 77.955 72.760 ;
        RECT 78.880 72.570 79.230 74.790 ;
        RECT 83.360 72.200 83.610 128.260 ;
        RECT 93.060 127.975 94.060 128.010 ;
        RECT 94.940 127.975 95.940 128.010 ;
        RECT 96.820 127.975 97.820 128.010 ;
        RECT 85.550 127.930 86.540 127.970 ;
        RECT 87.420 127.930 88.400 127.970 ;
        RECT 85.550 127.680 88.400 127.930 ;
        RECT 93.060 127.725 97.820 127.975 ;
        RECT 93.060 127.690 94.060 127.725 ;
        RECT 94.940 127.690 95.940 127.725 ;
        RECT 96.820 127.690 97.820 127.725 ;
        RECT 85.550 127.650 86.540 127.680 ;
        RECT 87.420 127.650 88.400 127.680 ;
        RECT 98.550 126.625 99.550 126.740 ;
        RECT 88.885 126.375 99.550 126.625 ;
        RECT 85.560 125.110 86.520 125.370 ;
        RECT 87.440 125.110 88.410 125.370 ;
        RECT 85.560 124.860 88.410 125.110 ;
        RECT 85.560 124.600 86.520 124.860 ;
        RECT 87.440 124.590 88.410 124.860 ;
        RECT 88.885 124.205 89.135 126.375 ;
        RECT 89.680 125.940 98.350 126.180 ;
        RECT 89.680 125.370 89.920 125.940 ;
        RECT 90.465 125.520 92.740 125.760 ;
        RECT 89.320 124.600 90.280 125.370 ;
        RECT 88.885 123.955 89.370 124.205 ;
        RECT 89.120 123.050 89.370 123.955 ;
        RECT 85.140 122.440 85.740 123.050 ;
        RECT 88.940 122.450 89.550 123.050 ;
        RECT 85.310 122.015 85.560 122.440 ;
        RECT 89.120 122.015 89.370 122.450 ;
        RECT 85.310 121.765 89.370 122.015 ;
        RECT 85.310 121.280 85.560 121.765 ;
        RECT 89.120 121.280 89.370 121.765 ;
        RECT 83.910 120.280 85.910 121.280 ;
        RECT 88.940 120.680 89.550 121.280 ;
        RECT 89.690 120.030 89.930 124.600 ;
        RECT 90.465 124.200 91.025 125.520 ;
        RECT 91.200 124.600 92.160 125.370 ;
        RECT 85.920 119.790 89.930 120.030 ;
        RECT 91.570 122.020 91.810 124.600 ;
        RECT 92.500 122.860 92.740 125.520 ;
        RECT 93.060 125.110 94.060 125.370 ;
        RECT 94.940 125.110 95.940 125.370 ;
        RECT 96.820 125.110 97.820 125.370 ;
        RECT 93.060 124.860 97.820 125.110 ;
        RECT 98.110 125.220 98.350 125.940 ;
        RECT 98.550 125.740 99.550 126.375 ;
        RECT 98.550 125.220 99.550 125.440 ;
        RECT 98.110 124.980 99.550 125.220 ;
        RECT 93.060 124.600 94.060 124.860 ;
        RECT 94.940 124.600 95.940 124.860 ;
        RECT 96.820 124.600 97.820 124.860 ;
        RECT 98.550 124.440 99.550 124.980 ;
        RECT 98.550 123.785 99.550 124.160 ;
        RECT 99.890 123.785 100.140 128.010 ;
        RECT 101.590 126.810 101.840 128.310 ;
        RECT 100.360 124.780 100.620 125.100 ;
        RECT 98.550 123.670 100.140 123.785 ;
        RECT 94.750 123.535 100.140 123.670 ;
        RECT 94.750 123.430 99.550 123.535 ;
        RECT 93.910 122.860 94.510 123.050 ;
        RECT 92.500 122.620 94.510 122.860 ;
        RECT 93.910 122.450 94.510 122.620 ;
        RECT 94.750 122.020 94.990 123.430 ;
        RECT 98.550 123.160 99.550 123.430 ;
        RECT 95.790 122.450 96.390 123.050 ;
        RECT 91.570 121.780 94.990 122.020 ;
        RECT 85.920 117.080 86.160 119.790 ;
        RECT 91.570 118.980 91.810 121.780 ;
        RECT 95.965 121.350 96.215 122.450 ;
        RECT 93.900 121.170 94.510 121.350 ;
        RECT 87.800 118.740 91.810 118.980 ;
        RECT 92.540 120.930 94.510 121.170 ;
        RECT 85.560 116.320 86.520 117.080 ;
        RECT 86.730 115.880 87.260 117.520 ;
        RECT 87.800 117.080 88.040 118.740 ;
        RECT 87.450 116.320 88.390 117.080 ;
        RECT 89.320 116.825 90.280 117.090 ;
        RECT 91.200 116.825 92.160 117.090 ;
        RECT 89.320 116.575 92.160 116.825 ;
        RECT 89.320 116.310 90.280 116.575 ;
        RECT 91.200 116.310 92.160 116.575 ;
        RECT 86.875 115.600 87.115 115.880 ;
        RECT 92.540 115.600 92.780 120.930 ;
        RECT 93.900 120.750 94.510 120.930 ;
        RECT 95.780 120.750 96.390 121.350 ;
        RECT 93.060 116.825 94.060 117.090 ;
        RECT 94.940 116.825 95.940 117.090 ;
        RECT 93.060 116.575 95.940 116.825 ;
        RECT 93.060 116.310 94.060 116.575 ;
        RECT 94.940 116.310 95.940 116.575 ;
        RECT 86.875 115.360 92.780 115.600 ;
        RECT 89.320 111.580 92.160 111.900 ;
        RECT 93.060 110.635 94.060 110.670 ;
        RECT 94.940 110.635 95.940 110.670 ;
        RECT 96.820 110.635 97.820 110.670 ;
        RECT 85.550 110.590 86.540 110.630 ;
        RECT 87.420 110.590 88.400 110.630 ;
        RECT 85.550 110.340 88.400 110.590 ;
        RECT 93.060 110.385 97.820 110.635 ;
        RECT 93.060 110.350 94.060 110.385 ;
        RECT 94.940 110.350 95.940 110.385 ;
        RECT 96.820 110.350 97.820 110.385 ;
        RECT 85.550 110.310 86.540 110.340 ;
        RECT 87.420 110.310 88.400 110.340 ;
        RECT 98.550 109.285 99.550 109.400 ;
        RECT 88.885 109.035 99.550 109.285 ;
        RECT 85.560 107.770 86.520 108.030 ;
        RECT 87.440 107.770 88.410 108.030 ;
        RECT 85.560 107.520 88.410 107.770 ;
        RECT 85.560 107.260 86.520 107.520 ;
        RECT 87.440 107.250 88.410 107.520 ;
        RECT 88.885 106.865 89.135 109.035 ;
        RECT 89.680 108.600 98.350 108.840 ;
        RECT 89.680 108.030 89.920 108.600 ;
        RECT 90.465 108.180 92.740 108.420 ;
        RECT 89.320 107.260 90.280 108.030 ;
        RECT 88.885 106.615 89.370 106.865 ;
        RECT 89.120 105.710 89.370 106.615 ;
        RECT 85.140 105.100 85.740 105.710 ;
        RECT 88.940 105.110 89.550 105.710 ;
        RECT 85.310 104.675 85.560 105.100 ;
        RECT 89.120 104.675 89.370 105.110 ;
        RECT 85.310 104.425 89.370 104.675 ;
        RECT 85.310 103.940 85.560 104.425 ;
        RECT 89.120 103.940 89.370 104.425 ;
        RECT 83.910 102.940 85.910 103.940 ;
        RECT 88.940 103.340 89.550 103.940 ;
        RECT 89.690 102.690 89.930 107.260 ;
        RECT 90.465 106.860 91.025 108.180 ;
        RECT 91.200 107.260 92.160 108.030 ;
        RECT 85.920 102.450 89.930 102.690 ;
        RECT 91.570 104.680 91.810 107.260 ;
        RECT 92.500 105.520 92.740 108.180 ;
        RECT 93.060 107.770 94.060 108.030 ;
        RECT 94.940 107.770 95.940 108.030 ;
        RECT 96.820 107.770 97.820 108.030 ;
        RECT 93.060 107.520 97.820 107.770 ;
        RECT 98.110 107.880 98.350 108.600 ;
        RECT 98.550 108.400 99.550 109.035 ;
        RECT 98.550 107.880 99.550 108.100 ;
        RECT 98.110 107.640 99.550 107.880 ;
        RECT 93.060 107.260 94.060 107.520 ;
        RECT 94.940 107.260 95.940 107.520 ;
        RECT 96.820 107.260 97.820 107.520 ;
        RECT 98.550 107.100 99.550 107.640 ;
        RECT 98.550 106.445 99.550 106.820 ;
        RECT 99.890 106.445 100.140 123.535 ;
        RECT 100.365 119.675 100.615 124.780 ;
        RECT 101.540 124.590 101.890 126.810 ;
        RECT 101.540 120.090 101.890 122.310 ;
        RECT 102.820 120.280 103.820 121.280 ;
        RECT 101.590 119.675 101.840 120.090 ;
        RECT 100.365 119.425 101.840 119.675 ;
        RECT 101.590 119.020 101.840 119.425 ;
        RECT 101.540 116.800 101.890 119.020 ;
        RECT 101.540 112.300 101.890 114.520 ;
        RECT 101.590 109.470 101.840 112.300 ;
        RECT 100.360 107.440 100.620 107.760 ;
        RECT 98.550 106.330 100.140 106.445 ;
        RECT 94.750 106.195 100.140 106.330 ;
        RECT 94.750 106.090 99.550 106.195 ;
        RECT 93.910 105.520 94.510 105.710 ;
        RECT 92.500 105.280 94.510 105.520 ;
        RECT 93.910 105.110 94.510 105.280 ;
        RECT 94.750 104.680 94.990 106.090 ;
        RECT 98.550 105.820 99.550 106.090 ;
        RECT 95.790 105.110 96.390 105.710 ;
        RECT 91.570 104.440 94.990 104.680 ;
        RECT 85.920 99.740 86.160 102.450 ;
        RECT 91.570 101.640 91.810 104.440 ;
        RECT 95.965 104.010 96.215 105.110 ;
        RECT 93.900 103.830 94.510 104.010 ;
        RECT 87.800 101.400 91.810 101.640 ;
        RECT 92.540 103.590 94.510 103.830 ;
        RECT 85.560 98.980 86.520 99.740 ;
        RECT 86.730 98.540 87.260 100.180 ;
        RECT 87.800 99.740 88.040 101.400 ;
        RECT 87.450 98.980 88.390 99.740 ;
        RECT 89.320 99.485 90.280 99.750 ;
        RECT 91.200 99.485 92.160 99.750 ;
        RECT 89.320 99.235 92.160 99.485 ;
        RECT 89.320 98.970 90.280 99.235 ;
        RECT 91.200 98.970 92.160 99.235 ;
        RECT 86.875 98.260 87.115 98.540 ;
        RECT 92.540 98.260 92.780 103.590 ;
        RECT 93.900 103.410 94.510 103.590 ;
        RECT 95.780 103.410 96.390 104.010 ;
        RECT 93.060 99.485 94.060 99.750 ;
        RECT 94.940 99.485 95.940 99.750 ;
        RECT 93.060 99.235 95.940 99.485 ;
        RECT 93.060 98.970 94.060 99.235 ;
        RECT 94.940 98.970 95.940 99.235 ;
        RECT 86.875 98.020 92.780 98.260 ;
        RECT 89.320 94.240 92.160 94.560 ;
        RECT 93.060 93.295 94.060 93.330 ;
        RECT 94.940 93.295 95.940 93.330 ;
        RECT 96.820 93.295 97.820 93.330 ;
        RECT 85.550 93.250 86.540 93.290 ;
        RECT 87.420 93.250 88.400 93.290 ;
        RECT 85.550 93.000 88.400 93.250 ;
        RECT 93.060 93.045 97.820 93.295 ;
        RECT 93.060 93.010 94.060 93.045 ;
        RECT 94.940 93.010 95.940 93.045 ;
        RECT 96.820 93.010 97.820 93.045 ;
        RECT 85.550 92.970 86.540 93.000 ;
        RECT 87.420 92.970 88.400 93.000 ;
        RECT 98.550 91.945 99.550 92.060 ;
        RECT 88.885 91.695 99.550 91.945 ;
        RECT 85.560 90.430 86.520 90.690 ;
        RECT 87.440 90.430 88.410 90.690 ;
        RECT 85.560 90.180 88.410 90.430 ;
        RECT 85.560 89.920 86.520 90.180 ;
        RECT 87.440 89.910 88.410 90.180 ;
        RECT 88.885 89.525 89.135 91.695 ;
        RECT 89.680 91.260 98.350 91.500 ;
        RECT 89.680 90.690 89.920 91.260 ;
        RECT 90.465 90.840 92.740 91.080 ;
        RECT 89.320 89.920 90.280 90.690 ;
        RECT 88.885 89.275 89.370 89.525 ;
        RECT 89.120 88.370 89.370 89.275 ;
        RECT 85.140 87.760 85.740 88.370 ;
        RECT 88.940 87.770 89.550 88.370 ;
        RECT 85.310 87.335 85.560 87.760 ;
        RECT 89.120 87.335 89.370 87.770 ;
        RECT 85.310 87.085 89.370 87.335 ;
        RECT 85.310 86.600 85.560 87.085 ;
        RECT 89.120 86.600 89.370 87.085 ;
        RECT 83.910 85.600 85.910 86.600 ;
        RECT 88.940 86.000 89.550 86.600 ;
        RECT 89.690 85.350 89.930 89.920 ;
        RECT 90.465 89.520 91.025 90.840 ;
        RECT 91.200 89.920 92.160 90.690 ;
        RECT 85.920 85.110 89.930 85.350 ;
        RECT 91.570 87.340 91.810 89.920 ;
        RECT 92.500 88.180 92.740 90.840 ;
        RECT 93.060 90.430 94.060 90.690 ;
        RECT 94.940 90.430 95.940 90.690 ;
        RECT 96.820 90.430 97.820 90.690 ;
        RECT 93.060 90.180 97.820 90.430 ;
        RECT 98.110 90.540 98.350 91.260 ;
        RECT 98.550 91.060 99.550 91.695 ;
        RECT 98.550 90.540 99.550 90.760 ;
        RECT 98.110 90.300 99.550 90.540 ;
        RECT 93.060 89.920 94.060 90.180 ;
        RECT 94.940 89.920 95.940 90.180 ;
        RECT 96.820 89.920 97.820 90.180 ;
        RECT 98.550 89.760 99.550 90.300 ;
        RECT 98.550 89.105 99.550 89.480 ;
        RECT 99.890 89.105 100.140 106.195 ;
        RECT 100.365 102.335 100.615 107.440 ;
        RECT 101.540 107.250 101.890 109.470 ;
        RECT 101.540 102.750 101.890 104.970 ;
        RECT 102.820 102.940 103.820 103.940 ;
        RECT 101.590 102.335 101.840 102.750 ;
        RECT 100.365 102.085 101.840 102.335 ;
        RECT 101.590 101.680 101.840 102.085 ;
        RECT 101.540 99.460 101.890 101.680 ;
        RECT 101.540 94.960 101.890 97.180 ;
        RECT 101.590 92.130 101.840 94.960 ;
        RECT 100.360 90.100 100.620 90.420 ;
        RECT 98.550 88.990 100.140 89.105 ;
        RECT 94.750 88.855 100.140 88.990 ;
        RECT 94.750 88.750 99.550 88.855 ;
        RECT 93.910 88.180 94.510 88.370 ;
        RECT 92.500 87.940 94.510 88.180 ;
        RECT 93.910 87.770 94.510 87.940 ;
        RECT 94.750 87.340 94.990 88.750 ;
        RECT 98.550 88.480 99.550 88.750 ;
        RECT 95.790 87.770 96.390 88.370 ;
        RECT 91.570 87.100 94.990 87.340 ;
        RECT 85.920 82.400 86.160 85.110 ;
        RECT 91.570 84.300 91.810 87.100 ;
        RECT 95.965 86.670 96.215 87.770 ;
        RECT 93.900 86.490 94.510 86.670 ;
        RECT 87.800 84.060 91.810 84.300 ;
        RECT 92.540 86.250 94.510 86.490 ;
        RECT 85.560 81.640 86.520 82.400 ;
        RECT 86.730 81.200 87.260 82.840 ;
        RECT 87.800 82.400 88.040 84.060 ;
        RECT 87.450 81.640 88.390 82.400 ;
        RECT 89.320 82.145 90.280 82.410 ;
        RECT 91.200 82.145 92.160 82.410 ;
        RECT 89.320 81.895 92.160 82.145 ;
        RECT 89.320 81.630 90.280 81.895 ;
        RECT 91.200 81.630 92.160 81.895 ;
        RECT 86.875 80.920 87.115 81.200 ;
        RECT 92.540 80.920 92.780 86.250 ;
        RECT 93.900 86.070 94.510 86.250 ;
        RECT 95.780 86.070 96.390 86.670 ;
        RECT 93.060 82.145 94.060 82.410 ;
        RECT 94.940 82.145 95.940 82.410 ;
        RECT 93.060 81.895 95.940 82.145 ;
        RECT 93.060 81.630 94.060 81.895 ;
        RECT 94.940 81.630 95.940 81.895 ;
        RECT 86.875 80.680 92.780 80.920 ;
        RECT 89.320 76.900 92.160 77.220 ;
        RECT 93.060 75.955 94.060 75.990 ;
        RECT 94.940 75.955 95.940 75.990 ;
        RECT 96.820 75.955 97.820 75.990 ;
        RECT 85.550 75.910 86.540 75.950 ;
        RECT 87.420 75.910 88.400 75.950 ;
        RECT 85.550 75.660 88.400 75.910 ;
        RECT 93.060 75.705 97.820 75.955 ;
        RECT 93.060 75.670 94.060 75.705 ;
        RECT 94.940 75.670 95.940 75.705 ;
        RECT 96.820 75.670 97.820 75.705 ;
        RECT 85.550 75.630 86.540 75.660 ;
        RECT 87.420 75.630 88.400 75.660 ;
        RECT 98.550 74.605 99.550 74.720 ;
        RECT 88.885 74.355 99.550 74.605 ;
        RECT 85.560 73.090 86.520 73.350 ;
        RECT 87.440 73.090 88.410 73.350 ;
        RECT 85.560 72.840 88.410 73.090 ;
        RECT 85.560 72.580 86.520 72.840 ;
        RECT 87.440 72.570 88.410 72.840 ;
        RECT 83.320 71.140 83.650 72.200 ;
        RECT 88.885 72.185 89.135 74.355 ;
        RECT 89.680 73.920 98.350 74.160 ;
        RECT 89.680 73.350 89.920 73.920 ;
        RECT 90.465 73.500 92.740 73.740 ;
        RECT 89.320 72.580 90.280 73.350 ;
        RECT 88.885 71.935 89.370 72.185 ;
        RECT 89.120 71.030 89.370 71.935 ;
        RECT 85.140 70.420 85.740 71.030 ;
        RECT 88.940 70.430 89.550 71.030 ;
        RECT 78.880 68.070 79.230 70.290 ;
        RECT 85.310 69.995 85.560 70.420 ;
        RECT 89.120 69.995 89.370 70.430 ;
        RECT 85.310 69.745 89.370 69.995 ;
        RECT 85.310 69.260 85.560 69.745 ;
        RECT 89.120 69.260 89.370 69.745 ;
        RECT 80.160 68.260 81.160 69.260 ;
        RECT 83.910 68.260 85.910 69.260 ;
        RECT 88.940 68.660 89.550 69.260 ;
        RECT 78.930 67.655 79.180 68.070 ;
        RECT 89.690 68.010 89.930 72.580 ;
        RECT 90.465 72.180 91.025 73.500 ;
        RECT 91.200 72.580 92.160 73.350 ;
        RECT 77.705 67.405 79.180 67.655 ;
        RECT 78.930 67.000 79.180 67.405 ;
        RECT 85.920 67.770 89.930 68.010 ;
        RECT 91.570 70.000 91.810 72.580 ;
        RECT 92.500 70.840 92.740 73.500 ;
        RECT 93.060 73.090 94.060 73.350 ;
        RECT 94.940 73.090 95.940 73.350 ;
        RECT 96.820 73.090 97.820 73.350 ;
        RECT 93.060 72.840 97.820 73.090 ;
        RECT 98.110 73.200 98.350 73.920 ;
        RECT 98.550 73.720 99.550 74.355 ;
        RECT 98.550 73.200 99.550 73.420 ;
        RECT 98.110 72.960 99.550 73.200 ;
        RECT 93.060 72.580 94.060 72.840 ;
        RECT 94.940 72.580 95.940 72.840 ;
        RECT 96.820 72.580 97.820 72.840 ;
        RECT 98.550 72.420 99.550 72.960 ;
        RECT 98.550 71.765 99.550 72.140 ;
        RECT 99.890 71.765 100.140 88.855 ;
        RECT 100.365 84.995 100.615 90.100 ;
        RECT 101.540 89.910 101.890 92.130 ;
        RECT 101.540 85.410 101.890 87.630 ;
        RECT 102.820 85.600 103.820 86.600 ;
        RECT 101.590 84.995 101.840 85.410 ;
        RECT 100.365 84.745 101.840 84.995 ;
        RECT 101.590 84.340 101.840 84.745 ;
        RECT 101.540 82.120 101.890 84.340 ;
        RECT 101.540 77.620 101.890 79.840 ;
        RECT 101.590 74.790 101.840 77.620 ;
        RECT 100.360 72.760 100.620 73.080 ;
        RECT 98.550 71.650 100.140 71.765 ;
        RECT 94.750 71.515 100.140 71.650 ;
        RECT 94.750 71.410 99.550 71.515 ;
        RECT 93.910 70.840 94.510 71.030 ;
        RECT 92.500 70.600 94.510 70.840 ;
        RECT 93.910 70.430 94.510 70.600 ;
        RECT 94.750 70.000 94.990 71.410 ;
        RECT 98.550 71.140 99.550 71.410 ;
        RECT 95.790 70.430 96.390 71.030 ;
        RECT 91.570 69.760 94.990 70.000 ;
        RECT 78.880 64.780 79.230 67.000 ;
        RECT 85.920 65.060 86.160 67.770 ;
        RECT 91.570 66.960 91.810 69.760 ;
        RECT 95.965 69.330 96.215 70.430 ;
        RECT 93.900 69.150 94.510 69.330 ;
        RECT 87.800 66.720 91.810 66.960 ;
        RECT 92.540 68.910 94.510 69.150 ;
        RECT 85.560 64.300 86.520 65.060 ;
        RECT 86.730 63.860 87.260 65.500 ;
        RECT 87.800 65.060 88.040 66.720 ;
        RECT 87.450 64.300 88.390 65.060 ;
        RECT 89.320 64.805 90.280 65.070 ;
        RECT 91.200 64.805 92.160 65.070 ;
        RECT 89.320 64.555 92.160 64.805 ;
        RECT 89.320 64.290 90.280 64.555 ;
        RECT 91.200 64.290 92.160 64.555 ;
        RECT 86.875 63.580 87.115 63.860 ;
        RECT 92.540 63.580 92.780 68.910 ;
        RECT 93.900 68.730 94.510 68.910 ;
        RECT 95.780 68.730 96.390 69.330 ;
        RECT 93.060 64.805 94.060 65.070 ;
        RECT 94.940 64.805 95.940 65.070 ;
        RECT 93.060 64.555 95.940 64.805 ;
        RECT 93.060 64.290 94.060 64.555 ;
        RECT 94.940 64.290 95.940 64.555 ;
        RECT 86.875 63.340 92.780 63.580 ;
        RECT 78.880 60.280 79.230 62.500 ;
        RECT 56.265 58.910 56.520 59.465 ;
        RECT 77.225 59.005 77.480 59.465 ;
        RECT 78.930 59.505 79.180 60.280 ;
        RECT 89.320 59.560 92.160 59.880 ;
        RECT 56.260 58.590 56.530 58.910 ;
        RECT 77.225 58.455 77.475 59.005 ;
        RECT 78.930 58.910 79.185 59.505 ;
        RECT 78.920 58.590 79.200 58.910 ;
        RECT 99.890 58.455 100.140 71.515 ;
        RECT 100.365 67.655 100.615 72.760 ;
        RECT 101.540 72.570 101.890 74.790 ;
        RECT 104.220 72.200 104.470 129.880 ;
        RECT 105.820 129.510 106.070 129.880 ;
        RECT 104.820 129.260 106.070 129.510 ;
        RECT 104.825 128.010 105.075 129.260 ;
        RECT 107.420 129.010 107.670 129.880 ;
        RECT 104.820 127.545 105.075 128.010 ;
        RECT 105.420 128.760 107.670 129.010 ;
        RECT 104.820 89.540 105.070 127.545 ;
        RECT 105.420 106.880 105.670 128.760 ;
        RECT 109.020 128.510 109.270 129.880 ;
        RECT 106.020 128.260 109.270 128.510 ;
        RECT 106.020 124.220 106.270 128.260 ;
        RECT 115.720 127.975 116.720 128.010 ;
        RECT 117.600 127.975 118.600 128.010 ;
        RECT 119.480 127.975 120.480 128.010 ;
        RECT 108.210 127.930 109.200 127.970 ;
        RECT 110.080 127.930 111.060 127.970 ;
        RECT 108.210 127.680 111.060 127.930 ;
        RECT 115.720 127.725 120.480 127.975 ;
        RECT 115.720 127.690 116.720 127.725 ;
        RECT 117.600 127.690 118.600 127.725 ;
        RECT 119.480 127.690 120.480 127.725 ;
        RECT 108.210 127.650 109.200 127.680 ;
        RECT 110.080 127.650 111.060 127.680 ;
        RECT 121.210 126.625 122.210 126.740 ;
        RECT 111.545 126.375 122.210 126.625 ;
        RECT 108.220 125.110 109.180 125.370 ;
        RECT 110.100 125.110 111.070 125.370 ;
        RECT 108.220 124.860 111.070 125.110 ;
        RECT 108.220 124.600 109.180 124.860 ;
        RECT 110.100 124.590 111.070 124.860 ;
        RECT 105.980 123.160 106.310 124.220 ;
        RECT 111.545 124.205 111.795 126.375 ;
        RECT 112.340 125.940 121.010 126.180 ;
        RECT 112.340 125.370 112.580 125.940 ;
        RECT 113.125 125.520 115.400 125.760 ;
        RECT 111.980 124.600 112.940 125.370 ;
        RECT 111.545 123.955 112.030 124.205 ;
        RECT 111.780 123.050 112.030 123.955 ;
        RECT 107.800 122.440 108.400 123.050 ;
        RECT 111.600 122.450 112.210 123.050 ;
        RECT 107.970 122.015 108.220 122.440 ;
        RECT 111.780 122.015 112.030 122.450 ;
        RECT 107.970 121.765 112.030 122.015 ;
        RECT 107.970 121.280 108.220 121.765 ;
        RECT 111.780 121.280 112.030 121.765 ;
        RECT 106.570 120.280 108.570 121.280 ;
        RECT 111.600 120.680 112.210 121.280 ;
        RECT 112.350 120.030 112.590 124.600 ;
        RECT 113.125 124.200 113.685 125.520 ;
        RECT 113.860 124.600 114.820 125.370 ;
        RECT 108.580 119.790 112.590 120.030 ;
        RECT 114.230 122.020 114.470 124.600 ;
        RECT 115.160 122.860 115.400 125.520 ;
        RECT 115.720 125.110 116.720 125.370 ;
        RECT 117.600 125.110 118.600 125.370 ;
        RECT 119.480 125.110 120.480 125.370 ;
        RECT 115.720 124.860 120.480 125.110 ;
        RECT 120.770 125.220 121.010 125.940 ;
        RECT 121.210 125.740 122.210 126.375 ;
        RECT 121.210 125.220 122.210 125.440 ;
        RECT 120.770 124.980 122.210 125.220 ;
        RECT 115.720 124.600 116.720 124.860 ;
        RECT 117.600 124.600 118.600 124.860 ;
        RECT 119.480 124.600 120.480 124.860 ;
        RECT 121.210 124.440 122.210 124.980 ;
        RECT 121.210 123.785 122.210 124.160 ;
        RECT 122.550 123.785 122.800 128.010 ;
        RECT 123.020 124.780 123.280 125.100 ;
        RECT 121.210 123.670 122.800 123.785 ;
        RECT 117.410 123.535 122.800 123.670 ;
        RECT 117.410 123.430 122.210 123.535 ;
        RECT 116.570 122.860 117.170 123.050 ;
        RECT 115.160 122.620 117.170 122.860 ;
        RECT 116.570 122.450 117.170 122.620 ;
        RECT 117.410 122.020 117.650 123.430 ;
        RECT 121.210 123.160 122.210 123.430 ;
        RECT 118.450 122.450 119.050 123.050 ;
        RECT 114.230 121.780 117.650 122.020 ;
        RECT 108.580 117.080 108.820 119.790 ;
        RECT 114.230 118.980 114.470 121.780 ;
        RECT 118.625 121.350 118.875 122.450 ;
        RECT 116.560 121.170 117.170 121.350 ;
        RECT 110.460 118.740 114.470 118.980 ;
        RECT 115.200 120.930 117.170 121.170 ;
        RECT 108.220 116.320 109.180 117.080 ;
        RECT 109.390 115.880 109.920 117.520 ;
        RECT 110.460 117.080 110.700 118.740 ;
        RECT 110.110 116.320 111.050 117.080 ;
        RECT 111.980 116.825 112.940 117.090 ;
        RECT 113.860 116.825 114.820 117.090 ;
        RECT 111.980 116.575 114.820 116.825 ;
        RECT 111.980 116.310 112.940 116.575 ;
        RECT 113.860 116.310 114.820 116.575 ;
        RECT 109.535 115.600 109.775 115.880 ;
        RECT 115.200 115.600 115.440 120.930 ;
        RECT 116.560 120.750 117.170 120.930 ;
        RECT 118.440 120.750 119.050 121.350 ;
        RECT 115.720 116.825 116.720 117.090 ;
        RECT 117.600 116.825 118.600 117.090 ;
        RECT 115.720 116.575 118.600 116.825 ;
        RECT 115.720 116.310 116.720 116.575 ;
        RECT 117.600 116.310 118.600 116.575 ;
        RECT 109.535 115.360 115.440 115.600 ;
        RECT 111.980 111.580 114.820 111.900 ;
        RECT 115.720 110.635 116.720 110.670 ;
        RECT 117.600 110.635 118.600 110.670 ;
        RECT 119.480 110.635 120.480 110.670 ;
        RECT 108.210 110.590 109.200 110.630 ;
        RECT 110.080 110.590 111.060 110.630 ;
        RECT 108.210 110.340 111.060 110.590 ;
        RECT 115.720 110.385 120.480 110.635 ;
        RECT 115.720 110.350 116.720 110.385 ;
        RECT 117.600 110.350 118.600 110.385 ;
        RECT 119.480 110.350 120.480 110.385 ;
        RECT 108.210 110.310 109.200 110.340 ;
        RECT 110.080 110.310 111.060 110.340 ;
        RECT 121.210 109.285 122.210 109.400 ;
        RECT 111.545 109.035 122.210 109.285 ;
        RECT 108.220 107.770 109.180 108.030 ;
        RECT 110.100 107.770 111.070 108.030 ;
        RECT 108.220 107.520 111.070 107.770 ;
        RECT 108.220 107.260 109.180 107.520 ;
        RECT 110.100 107.250 111.070 107.520 ;
        RECT 105.380 105.820 105.710 106.880 ;
        RECT 111.545 106.865 111.795 109.035 ;
        RECT 112.340 108.600 121.010 108.840 ;
        RECT 112.340 108.030 112.580 108.600 ;
        RECT 113.125 108.180 115.400 108.420 ;
        RECT 111.980 107.260 112.940 108.030 ;
        RECT 111.545 106.615 112.030 106.865 ;
        RECT 111.780 105.710 112.030 106.615 ;
        RECT 107.800 105.100 108.400 105.710 ;
        RECT 111.600 105.110 112.210 105.710 ;
        RECT 107.970 104.675 108.220 105.100 ;
        RECT 111.780 104.675 112.030 105.110 ;
        RECT 107.970 104.425 112.030 104.675 ;
        RECT 107.970 103.940 108.220 104.425 ;
        RECT 111.780 103.940 112.030 104.425 ;
        RECT 106.570 102.940 108.570 103.940 ;
        RECT 111.600 103.340 112.210 103.940 ;
        RECT 112.350 102.690 112.590 107.260 ;
        RECT 113.125 106.860 113.685 108.180 ;
        RECT 113.860 107.260 114.820 108.030 ;
        RECT 108.580 102.450 112.590 102.690 ;
        RECT 114.230 104.680 114.470 107.260 ;
        RECT 115.160 105.520 115.400 108.180 ;
        RECT 115.720 107.770 116.720 108.030 ;
        RECT 117.600 107.770 118.600 108.030 ;
        RECT 119.480 107.770 120.480 108.030 ;
        RECT 115.720 107.520 120.480 107.770 ;
        RECT 120.770 107.880 121.010 108.600 ;
        RECT 121.210 108.400 122.210 109.035 ;
        RECT 121.210 107.880 122.210 108.100 ;
        RECT 120.770 107.640 122.210 107.880 ;
        RECT 115.720 107.260 116.720 107.520 ;
        RECT 117.600 107.260 118.600 107.520 ;
        RECT 119.480 107.260 120.480 107.520 ;
        RECT 121.210 107.100 122.210 107.640 ;
        RECT 121.210 106.445 122.210 106.820 ;
        RECT 122.550 106.445 122.800 123.535 ;
        RECT 123.025 119.675 123.275 124.780 ;
        RECT 124.200 120.090 124.550 122.310 ;
        RECT 124.250 119.675 124.500 120.090 ;
        RECT 123.025 119.425 124.500 119.675 ;
        RECT 124.250 119.020 124.500 119.425 ;
        RECT 124.200 116.800 124.550 119.020 ;
        RECT 124.200 112.300 124.550 114.520 ;
        RECT 124.250 109.470 124.500 112.300 ;
        RECT 123.020 107.440 123.280 107.760 ;
        RECT 121.210 106.330 122.800 106.445 ;
        RECT 117.410 106.195 122.800 106.330 ;
        RECT 117.410 106.090 122.210 106.195 ;
        RECT 116.570 105.520 117.170 105.710 ;
        RECT 115.160 105.280 117.170 105.520 ;
        RECT 116.570 105.110 117.170 105.280 ;
        RECT 117.410 104.680 117.650 106.090 ;
        RECT 121.210 105.820 122.210 106.090 ;
        RECT 118.450 105.110 119.050 105.710 ;
        RECT 114.230 104.440 117.650 104.680 ;
        RECT 108.580 99.740 108.820 102.450 ;
        RECT 114.230 101.640 114.470 104.440 ;
        RECT 118.625 104.010 118.875 105.110 ;
        RECT 116.560 103.830 117.170 104.010 ;
        RECT 110.460 101.400 114.470 101.640 ;
        RECT 115.200 103.590 117.170 103.830 ;
        RECT 108.220 98.980 109.180 99.740 ;
        RECT 109.390 98.540 109.920 100.180 ;
        RECT 110.460 99.740 110.700 101.400 ;
        RECT 110.110 98.980 111.050 99.740 ;
        RECT 111.980 99.485 112.940 99.750 ;
        RECT 113.860 99.485 114.820 99.750 ;
        RECT 111.980 99.235 114.820 99.485 ;
        RECT 111.980 98.970 112.940 99.235 ;
        RECT 113.860 98.970 114.820 99.235 ;
        RECT 109.535 98.260 109.775 98.540 ;
        RECT 115.200 98.260 115.440 103.590 ;
        RECT 116.560 103.410 117.170 103.590 ;
        RECT 118.440 103.410 119.050 104.010 ;
        RECT 115.720 99.485 116.720 99.750 ;
        RECT 117.600 99.485 118.600 99.750 ;
        RECT 115.720 99.235 118.600 99.485 ;
        RECT 115.720 98.970 116.720 99.235 ;
        RECT 117.600 98.970 118.600 99.235 ;
        RECT 109.535 98.020 115.440 98.260 ;
        RECT 111.980 94.240 114.820 94.560 ;
        RECT 115.720 93.295 116.720 93.330 ;
        RECT 117.600 93.295 118.600 93.330 ;
        RECT 119.480 93.295 120.480 93.330 ;
        RECT 108.210 93.250 109.200 93.290 ;
        RECT 110.080 93.250 111.060 93.290 ;
        RECT 108.210 93.000 111.060 93.250 ;
        RECT 115.720 93.045 120.480 93.295 ;
        RECT 115.720 93.010 116.720 93.045 ;
        RECT 117.600 93.010 118.600 93.045 ;
        RECT 119.480 93.010 120.480 93.045 ;
        RECT 108.210 92.970 109.200 93.000 ;
        RECT 110.080 92.970 111.060 93.000 ;
        RECT 121.210 91.945 122.210 92.060 ;
        RECT 111.545 91.695 122.210 91.945 ;
        RECT 108.220 90.430 109.180 90.690 ;
        RECT 110.100 90.430 111.070 90.690 ;
        RECT 108.220 90.180 111.070 90.430 ;
        RECT 108.220 89.920 109.180 90.180 ;
        RECT 110.100 89.910 111.070 90.180 ;
        RECT 104.780 88.480 105.110 89.540 ;
        RECT 111.545 89.525 111.795 91.695 ;
        RECT 112.340 91.260 121.010 91.500 ;
        RECT 112.340 90.690 112.580 91.260 ;
        RECT 113.125 90.840 115.400 91.080 ;
        RECT 111.980 89.920 112.940 90.690 ;
        RECT 111.545 89.275 112.030 89.525 ;
        RECT 111.780 88.370 112.030 89.275 ;
        RECT 107.800 87.760 108.400 88.370 ;
        RECT 111.600 87.770 112.210 88.370 ;
        RECT 107.970 87.335 108.220 87.760 ;
        RECT 111.780 87.335 112.030 87.770 ;
        RECT 107.970 87.085 112.030 87.335 ;
        RECT 107.970 86.600 108.220 87.085 ;
        RECT 111.780 86.600 112.030 87.085 ;
        RECT 106.570 85.600 108.570 86.600 ;
        RECT 111.600 86.000 112.210 86.600 ;
        RECT 112.350 85.350 112.590 89.920 ;
        RECT 113.125 89.520 113.685 90.840 ;
        RECT 113.860 89.920 114.820 90.690 ;
        RECT 108.580 85.110 112.590 85.350 ;
        RECT 114.230 87.340 114.470 89.920 ;
        RECT 115.160 88.180 115.400 90.840 ;
        RECT 115.720 90.430 116.720 90.690 ;
        RECT 117.600 90.430 118.600 90.690 ;
        RECT 119.480 90.430 120.480 90.690 ;
        RECT 115.720 90.180 120.480 90.430 ;
        RECT 120.770 90.540 121.010 91.260 ;
        RECT 121.210 91.060 122.210 91.695 ;
        RECT 121.210 90.540 122.210 90.760 ;
        RECT 120.770 90.300 122.210 90.540 ;
        RECT 115.720 89.920 116.720 90.180 ;
        RECT 117.600 89.920 118.600 90.180 ;
        RECT 119.480 89.920 120.480 90.180 ;
        RECT 121.210 89.760 122.210 90.300 ;
        RECT 121.210 89.105 122.210 89.480 ;
        RECT 122.550 89.105 122.800 106.195 ;
        RECT 123.025 102.335 123.275 107.440 ;
        RECT 124.200 107.250 124.550 109.470 ;
        RECT 124.200 102.750 124.550 104.970 ;
        RECT 124.250 102.335 124.500 102.750 ;
        RECT 123.025 102.085 124.500 102.335 ;
        RECT 124.250 101.680 124.500 102.085 ;
        RECT 124.200 99.460 124.550 101.680 ;
        RECT 124.200 94.960 124.550 97.180 ;
        RECT 124.250 92.130 124.500 94.960 ;
        RECT 123.020 90.100 123.280 90.420 ;
        RECT 121.210 88.990 122.800 89.105 ;
        RECT 117.410 88.855 122.800 88.990 ;
        RECT 117.410 88.750 122.210 88.855 ;
        RECT 116.570 88.180 117.170 88.370 ;
        RECT 115.160 87.940 117.170 88.180 ;
        RECT 116.570 87.770 117.170 87.940 ;
        RECT 117.410 87.340 117.650 88.750 ;
        RECT 121.210 88.480 122.210 88.750 ;
        RECT 118.450 87.770 119.050 88.370 ;
        RECT 114.230 87.100 117.650 87.340 ;
        RECT 108.580 82.400 108.820 85.110 ;
        RECT 114.230 84.300 114.470 87.100 ;
        RECT 118.625 86.670 118.875 87.770 ;
        RECT 116.560 86.490 117.170 86.670 ;
        RECT 110.460 84.060 114.470 84.300 ;
        RECT 115.200 86.250 117.170 86.490 ;
        RECT 108.220 81.640 109.180 82.400 ;
        RECT 109.390 81.200 109.920 82.840 ;
        RECT 110.460 82.400 110.700 84.060 ;
        RECT 110.110 81.640 111.050 82.400 ;
        RECT 111.980 82.145 112.940 82.410 ;
        RECT 113.860 82.145 114.820 82.410 ;
        RECT 111.980 81.895 114.820 82.145 ;
        RECT 111.980 81.630 112.940 81.895 ;
        RECT 113.860 81.630 114.820 81.895 ;
        RECT 109.535 80.920 109.775 81.200 ;
        RECT 115.200 80.920 115.440 86.250 ;
        RECT 116.560 86.070 117.170 86.250 ;
        RECT 118.440 86.070 119.050 86.670 ;
        RECT 115.720 82.145 116.720 82.410 ;
        RECT 117.600 82.145 118.600 82.410 ;
        RECT 115.720 81.895 118.600 82.145 ;
        RECT 115.720 81.630 116.720 81.895 ;
        RECT 117.600 81.630 118.600 81.895 ;
        RECT 109.535 80.680 115.440 80.920 ;
        RECT 111.980 76.900 114.820 77.220 ;
        RECT 115.720 75.955 116.720 75.990 ;
        RECT 117.600 75.955 118.600 75.990 ;
        RECT 119.480 75.955 120.480 75.990 ;
        RECT 108.210 75.910 109.200 75.950 ;
        RECT 110.080 75.910 111.060 75.950 ;
        RECT 108.210 75.660 111.060 75.910 ;
        RECT 115.720 75.705 120.480 75.955 ;
        RECT 115.720 75.670 116.720 75.705 ;
        RECT 117.600 75.670 118.600 75.705 ;
        RECT 119.480 75.670 120.480 75.705 ;
        RECT 108.210 75.630 109.200 75.660 ;
        RECT 110.080 75.630 111.060 75.660 ;
        RECT 121.210 74.605 122.210 74.720 ;
        RECT 111.545 74.355 122.210 74.605 ;
        RECT 108.220 73.090 109.180 73.350 ;
        RECT 110.100 73.090 111.070 73.350 ;
        RECT 108.220 72.840 111.070 73.090 ;
        RECT 108.220 72.580 109.180 72.840 ;
        RECT 110.100 72.570 111.070 72.840 ;
        RECT 104.180 71.140 104.510 72.200 ;
        RECT 111.545 72.185 111.795 74.355 ;
        RECT 112.340 73.920 121.010 74.160 ;
        RECT 112.340 73.350 112.580 73.920 ;
        RECT 113.125 73.500 115.400 73.740 ;
        RECT 111.980 72.580 112.940 73.350 ;
        RECT 111.545 71.935 112.030 72.185 ;
        RECT 111.780 71.030 112.030 71.935 ;
        RECT 107.800 70.420 108.400 71.030 ;
        RECT 111.600 70.430 112.210 71.030 ;
        RECT 101.540 68.070 101.890 70.290 ;
        RECT 107.970 69.995 108.220 70.420 ;
        RECT 111.780 69.995 112.030 70.430 ;
        RECT 107.970 69.745 112.030 69.995 ;
        RECT 107.970 69.260 108.220 69.745 ;
        RECT 111.780 69.260 112.030 69.745 ;
        RECT 102.820 68.260 103.820 69.260 ;
        RECT 106.570 68.260 108.570 69.260 ;
        RECT 111.600 68.660 112.210 69.260 ;
        RECT 101.590 67.655 101.840 68.070 ;
        RECT 112.350 68.010 112.590 72.580 ;
        RECT 113.125 72.180 113.685 73.500 ;
        RECT 113.860 72.580 114.820 73.350 ;
        RECT 100.365 67.405 101.840 67.655 ;
        RECT 101.590 67.000 101.840 67.405 ;
        RECT 108.580 67.770 112.590 68.010 ;
        RECT 114.230 70.000 114.470 72.580 ;
        RECT 115.160 70.840 115.400 73.500 ;
        RECT 115.720 73.090 116.720 73.350 ;
        RECT 117.600 73.090 118.600 73.350 ;
        RECT 119.480 73.090 120.480 73.350 ;
        RECT 115.720 72.840 120.480 73.090 ;
        RECT 120.770 73.200 121.010 73.920 ;
        RECT 121.210 73.720 122.210 74.355 ;
        RECT 121.210 73.200 122.210 73.420 ;
        RECT 120.770 72.960 122.210 73.200 ;
        RECT 115.720 72.580 116.720 72.840 ;
        RECT 117.600 72.580 118.600 72.840 ;
        RECT 119.480 72.580 120.480 72.840 ;
        RECT 121.210 72.420 122.210 72.960 ;
        RECT 121.210 71.765 122.210 72.140 ;
        RECT 122.550 71.765 122.800 88.855 ;
        RECT 123.025 84.995 123.275 90.100 ;
        RECT 124.200 89.910 124.550 92.130 ;
        RECT 124.200 85.410 124.550 87.630 ;
        RECT 124.250 84.995 124.500 85.410 ;
        RECT 123.025 84.745 124.500 84.995 ;
        RECT 124.250 84.340 124.500 84.745 ;
        RECT 124.200 82.120 124.550 84.340 ;
        RECT 124.200 77.620 124.550 79.840 ;
        RECT 124.250 74.790 124.500 77.620 ;
        RECT 123.020 72.760 123.280 73.080 ;
        RECT 121.210 71.650 122.800 71.765 ;
        RECT 117.410 71.515 122.800 71.650 ;
        RECT 117.410 71.410 122.210 71.515 ;
        RECT 116.570 70.840 117.170 71.030 ;
        RECT 115.160 70.600 117.170 70.840 ;
        RECT 116.570 70.430 117.170 70.600 ;
        RECT 117.410 70.000 117.650 71.410 ;
        RECT 121.210 71.140 122.210 71.410 ;
        RECT 118.450 70.430 119.050 71.030 ;
        RECT 114.230 69.760 117.650 70.000 ;
        RECT 101.540 64.780 101.890 67.000 ;
        RECT 108.580 65.060 108.820 67.770 ;
        RECT 114.230 66.960 114.470 69.760 ;
        RECT 118.625 69.330 118.875 70.430 ;
        RECT 116.560 69.150 117.170 69.330 ;
        RECT 110.460 66.720 114.470 66.960 ;
        RECT 115.200 68.910 117.170 69.150 ;
        RECT 108.220 64.300 109.180 65.060 ;
        RECT 109.390 63.860 109.920 65.500 ;
        RECT 110.460 65.060 110.700 66.720 ;
        RECT 110.110 64.300 111.050 65.060 ;
        RECT 111.980 64.805 112.940 65.070 ;
        RECT 113.860 64.805 114.820 65.070 ;
        RECT 111.980 64.555 114.820 64.805 ;
        RECT 111.980 64.290 112.940 64.555 ;
        RECT 113.860 64.290 114.820 64.555 ;
        RECT 109.535 63.580 109.775 63.860 ;
        RECT 115.200 63.580 115.440 68.910 ;
        RECT 116.560 68.730 117.170 68.910 ;
        RECT 118.440 68.730 119.050 69.330 ;
        RECT 115.720 64.805 116.720 65.070 ;
        RECT 117.600 64.805 118.600 65.070 ;
        RECT 115.720 64.555 118.600 64.805 ;
        RECT 115.720 64.290 116.720 64.555 ;
        RECT 117.600 64.290 118.600 64.555 ;
        RECT 109.535 63.340 115.440 63.580 ;
        RECT 101.540 60.280 101.890 62.500 ;
        RECT 101.590 59.875 101.840 60.280 ;
        RECT 101.590 58.910 101.845 59.875 ;
        RECT 111.980 59.560 114.820 59.880 ;
        RECT 101.580 58.590 101.850 58.910 ;
        RECT 122.550 58.455 122.800 71.515 ;
        RECT 123.025 67.655 123.275 72.760 ;
        RECT 124.200 72.570 124.550 74.790 ;
        RECT 124.200 68.070 124.550 70.290 ;
        RECT 124.250 67.655 124.500 68.070 ;
        RECT 123.025 67.405 124.500 67.655 ;
        RECT 124.250 67.000 124.500 67.405 ;
        RECT 124.200 64.780 124.550 67.000 ;
        RECT 124.200 60.280 124.550 62.500 ;
        RECT 124.250 58.910 124.500 60.280 ;
        RECT 124.245 58.590 124.505 58.910 ;
        RECT 38.875 58.205 54.820 58.455 ;
        RECT 61.535 58.205 77.480 58.455 ;
        RECT 84.195 58.205 100.140 58.455 ;
        RECT 106.855 58.205 122.800 58.455 ;
        RECT 38.875 50.885 39.125 58.205 ;
        RECT 47.740 57.955 48.740 57.990 ;
        RECT 49.620 57.955 50.620 57.990 ;
        RECT 51.500 57.955 52.500 57.990 ;
        RECT 40.230 57.910 41.220 57.950 ;
        RECT 42.100 57.910 43.080 57.950 ;
        RECT 40.230 57.660 43.080 57.910 ;
        RECT 47.740 57.705 52.500 57.955 ;
        RECT 47.740 57.670 48.740 57.705 ;
        RECT 49.620 57.670 50.620 57.705 ;
        RECT 51.500 57.670 52.500 57.705 ;
        RECT 40.230 57.630 41.220 57.660 ;
        RECT 42.100 57.630 43.080 57.660 ;
        RECT 53.230 56.605 54.230 56.720 ;
        RECT 43.565 56.355 54.230 56.605 ;
        RECT 40.240 55.090 41.200 55.350 ;
        RECT 42.120 55.090 43.090 55.350 ;
        RECT 40.240 54.840 43.090 55.090 ;
        RECT 40.240 54.580 41.200 54.840 ;
        RECT 42.120 54.570 43.090 54.840 ;
        RECT 43.565 54.185 43.815 56.355 ;
        RECT 44.360 55.920 53.030 56.160 ;
        RECT 44.360 55.350 44.600 55.920 ;
        RECT 45.145 55.500 47.420 55.740 ;
        RECT 44.000 54.580 44.960 55.350 ;
        RECT 43.565 53.935 44.050 54.185 ;
        RECT 43.795 53.030 44.050 53.935 ;
        RECT 39.820 52.420 40.420 53.030 ;
        RECT 43.620 52.430 44.230 53.030 ;
        RECT 39.990 51.995 40.240 52.420 ;
        RECT 43.795 51.995 44.050 52.430 ;
        RECT 39.990 51.745 44.050 51.995 ;
        RECT 39.990 51.465 40.245 51.745 ;
        RECT 39.990 51.260 40.240 51.465 ;
        RECT 43.800 51.260 44.050 51.745 ;
        RECT 39.590 50.885 40.590 51.260 ;
        RECT 38.875 50.635 40.590 50.885 ;
        RECT 43.620 50.660 44.230 51.260 ;
        RECT 39.590 50.260 40.590 50.635 ;
        RECT 44.370 50.010 44.610 54.580 ;
        RECT 45.145 54.180 45.705 55.500 ;
        RECT 47.180 52.840 47.420 55.500 ;
        RECT 47.740 55.090 48.740 55.350 ;
        RECT 49.620 55.090 50.620 55.350 ;
        RECT 51.500 55.090 52.500 55.350 ;
        RECT 47.740 54.840 52.500 55.090 ;
        RECT 52.790 55.200 53.030 55.920 ;
        RECT 53.230 55.720 54.230 56.355 ;
        RECT 53.605 55.420 53.855 55.720 ;
        RECT 53.230 55.200 54.230 55.420 ;
        RECT 52.790 54.960 54.230 55.200 ;
        RECT 47.740 54.580 48.740 54.840 ;
        RECT 49.620 54.580 50.620 54.840 ;
        RECT 51.500 54.580 52.500 54.840 ;
        RECT 53.230 54.420 54.230 54.960 ;
        RECT 48.590 52.840 49.190 53.030 ;
        RECT 47.180 52.600 49.190 52.840 ;
        RECT 48.590 52.430 49.190 52.600 ;
        RECT 50.470 52.430 51.070 53.030 ;
        RECT 50.645 51.330 50.895 52.430 ;
        RECT 48.580 51.150 49.190 51.330 ;
        RECT 40.600 49.770 44.610 50.010 ;
        RECT 47.220 50.910 49.190 51.150 ;
        RECT 40.600 47.060 40.840 49.770 ;
        RECT 40.240 46.300 41.200 47.060 ;
        RECT 41.410 45.860 41.940 47.500 ;
        RECT 44.000 46.805 44.960 47.070 ;
        RECT 45.880 46.805 46.840 47.070 ;
        RECT 44.000 46.555 46.840 46.805 ;
        RECT 44.000 46.290 44.960 46.555 ;
        RECT 45.880 46.290 46.840 46.555 ;
        RECT 41.555 45.580 41.795 45.860 ;
        RECT 47.220 45.580 47.460 50.910 ;
        RECT 48.580 50.730 49.190 50.910 ;
        RECT 50.460 50.730 51.070 51.330 ;
        RECT 61.535 50.885 61.785 58.205 ;
        RECT 70.400 57.955 71.400 57.990 ;
        RECT 72.280 57.955 73.280 57.990 ;
        RECT 74.160 57.955 75.160 57.990 ;
        RECT 62.890 57.910 63.880 57.950 ;
        RECT 64.760 57.910 65.740 57.950 ;
        RECT 62.890 57.660 65.740 57.910 ;
        RECT 70.400 57.705 75.160 57.955 ;
        RECT 70.400 57.670 71.400 57.705 ;
        RECT 72.280 57.670 73.280 57.705 ;
        RECT 74.160 57.670 75.160 57.705 ;
        RECT 62.890 57.630 63.880 57.660 ;
        RECT 64.760 57.630 65.740 57.660 ;
        RECT 75.890 56.605 76.890 56.720 ;
        RECT 66.225 56.355 76.890 56.605 ;
        RECT 62.900 55.090 63.860 55.350 ;
        RECT 64.780 55.090 65.750 55.350 ;
        RECT 62.900 54.840 65.750 55.090 ;
        RECT 62.900 54.580 63.860 54.840 ;
        RECT 64.780 54.570 65.750 54.840 ;
        RECT 66.225 54.185 66.475 56.355 ;
        RECT 67.020 55.920 75.690 56.160 ;
        RECT 67.020 55.350 67.260 55.920 ;
        RECT 67.805 55.500 70.080 55.740 ;
        RECT 66.660 54.580 67.620 55.350 ;
        RECT 66.225 53.935 66.710 54.185 ;
        RECT 66.455 53.030 66.710 53.935 ;
        RECT 62.480 52.420 63.080 53.030 ;
        RECT 66.280 52.430 66.890 53.030 ;
        RECT 62.650 51.995 62.900 52.420 ;
        RECT 66.455 51.995 66.710 52.430 ;
        RECT 62.650 51.745 66.710 51.995 ;
        RECT 62.650 51.465 62.905 51.745 ;
        RECT 62.650 51.260 62.900 51.465 ;
        RECT 66.460 51.260 66.710 51.745 ;
        RECT 62.250 50.885 63.250 51.260 ;
        RECT 61.535 50.635 63.250 50.885 ;
        RECT 66.280 50.660 66.890 51.260 ;
        RECT 62.250 50.260 63.250 50.635 ;
        RECT 67.030 50.010 67.270 54.580 ;
        RECT 67.805 54.180 68.365 55.500 ;
        RECT 69.840 52.840 70.080 55.500 ;
        RECT 70.400 55.090 71.400 55.350 ;
        RECT 72.280 55.090 73.280 55.350 ;
        RECT 74.160 55.090 75.160 55.350 ;
        RECT 70.400 54.840 75.160 55.090 ;
        RECT 75.450 55.200 75.690 55.920 ;
        RECT 75.890 55.720 76.890 56.355 ;
        RECT 76.265 55.420 76.515 55.720 ;
        RECT 75.890 55.200 76.890 55.420 ;
        RECT 75.450 54.960 76.890 55.200 ;
        RECT 70.400 54.580 71.400 54.840 ;
        RECT 72.280 54.580 73.280 54.840 ;
        RECT 74.160 54.580 75.160 54.840 ;
        RECT 75.890 54.420 76.890 54.960 ;
        RECT 71.250 52.840 71.850 53.030 ;
        RECT 69.840 52.600 71.850 52.840 ;
        RECT 71.250 52.430 71.850 52.600 ;
        RECT 73.130 52.430 73.730 53.030 ;
        RECT 73.305 51.330 73.555 52.430 ;
        RECT 71.240 51.150 71.850 51.330 ;
        RECT 63.260 49.770 67.270 50.010 ;
        RECT 69.880 50.910 71.850 51.150 ;
        RECT 47.740 46.805 48.740 47.070 ;
        RECT 49.620 46.805 50.620 47.070 ;
        RECT 63.260 47.060 63.500 49.770 ;
        RECT 47.740 46.555 50.620 46.805 ;
        RECT 47.740 46.290 48.740 46.555 ;
        RECT 49.620 46.290 50.620 46.555 ;
        RECT 62.900 46.300 63.860 47.060 ;
        RECT 64.070 45.860 64.600 47.500 ;
        RECT 66.660 46.805 67.620 47.070 ;
        RECT 68.540 46.805 69.500 47.070 ;
        RECT 66.660 46.555 69.500 46.805 ;
        RECT 66.660 46.290 67.620 46.555 ;
        RECT 68.540 46.290 69.500 46.555 ;
        RECT 41.555 45.340 47.460 45.580 ;
        RECT 64.215 45.580 64.455 45.860 ;
        RECT 69.880 45.580 70.120 50.910 ;
        RECT 71.240 50.730 71.850 50.910 ;
        RECT 73.120 50.730 73.730 51.330 ;
        RECT 84.195 50.885 84.445 58.205 ;
        RECT 93.060 57.955 94.060 57.990 ;
        RECT 94.940 57.955 95.940 57.990 ;
        RECT 96.820 57.955 97.820 57.990 ;
        RECT 85.550 57.910 86.540 57.950 ;
        RECT 87.420 57.910 88.400 57.950 ;
        RECT 85.550 57.660 88.400 57.910 ;
        RECT 93.060 57.705 97.820 57.955 ;
        RECT 93.060 57.670 94.060 57.705 ;
        RECT 94.940 57.670 95.940 57.705 ;
        RECT 96.820 57.670 97.820 57.705 ;
        RECT 85.550 57.630 86.540 57.660 ;
        RECT 87.420 57.630 88.400 57.660 ;
        RECT 98.550 56.605 99.550 56.720 ;
        RECT 88.885 56.355 99.550 56.605 ;
        RECT 85.560 55.090 86.520 55.350 ;
        RECT 87.440 55.090 88.410 55.350 ;
        RECT 85.560 54.840 88.410 55.090 ;
        RECT 85.560 54.580 86.520 54.840 ;
        RECT 87.440 54.570 88.410 54.840 ;
        RECT 88.885 54.185 89.135 56.355 ;
        RECT 89.680 55.920 98.350 56.160 ;
        RECT 89.680 55.350 89.920 55.920 ;
        RECT 90.465 55.500 92.740 55.740 ;
        RECT 89.320 54.580 90.280 55.350 ;
        RECT 88.885 53.935 89.370 54.185 ;
        RECT 89.115 53.030 89.370 53.935 ;
        RECT 85.140 52.420 85.740 53.030 ;
        RECT 88.940 52.430 89.550 53.030 ;
        RECT 85.310 51.995 85.560 52.420 ;
        RECT 89.115 51.995 89.370 52.430 ;
        RECT 85.310 51.745 89.370 51.995 ;
        RECT 85.310 51.465 85.565 51.745 ;
        RECT 85.310 51.260 85.560 51.465 ;
        RECT 89.120 51.260 89.370 51.745 ;
        RECT 84.910 50.885 85.910 51.260 ;
        RECT 84.195 50.635 85.910 50.885 ;
        RECT 88.940 50.660 89.550 51.260 ;
        RECT 84.910 50.260 85.910 50.635 ;
        RECT 89.690 50.010 89.930 54.580 ;
        RECT 90.465 54.180 91.025 55.500 ;
        RECT 92.500 52.840 92.740 55.500 ;
        RECT 93.060 55.090 94.060 55.350 ;
        RECT 94.940 55.090 95.940 55.350 ;
        RECT 96.820 55.090 97.820 55.350 ;
        RECT 93.060 54.840 97.820 55.090 ;
        RECT 98.110 55.200 98.350 55.920 ;
        RECT 98.550 55.720 99.550 56.355 ;
        RECT 98.925 55.420 99.175 55.720 ;
        RECT 98.550 55.200 99.550 55.420 ;
        RECT 98.110 54.960 99.550 55.200 ;
        RECT 93.060 54.580 94.060 54.840 ;
        RECT 94.940 54.580 95.940 54.840 ;
        RECT 96.820 54.580 97.820 54.840 ;
        RECT 98.550 54.420 99.550 54.960 ;
        RECT 93.910 52.840 94.510 53.030 ;
        RECT 92.500 52.600 94.510 52.840 ;
        RECT 93.910 52.430 94.510 52.600 ;
        RECT 95.790 52.430 96.390 53.030 ;
        RECT 95.965 51.330 96.215 52.430 ;
        RECT 93.900 51.150 94.510 51.330 ;
        RECT 85.920 49.770 89.930 50.010 ;
        RECT 92.540 50.910 94.510 51.150 ;
        RECT 70.400 46.805 71.400 47.070 ;
        RECT 72.280 46.805 73.280 47.070 ;
        RECT 85.920 47.060 86.160 49.770 ;
        RECT 70.400 46.555 73.280 46.805 ;
        RECT 70.400 46.290 71.400 46.555 ;
        RECT 72.280 46.290 73.280 46.555 ;
        RECT 85.560 46.300 86.520 47.060 ;
        RECT 86.730 45.860 87.260 47.500 ;
        RECT 89.320 46.805 90.280 47.070 ;
        RECT 91.200 46.805 92.160 47.070 ;
        RECT 89.320 46.555 92.160 46.805 ;
        RECT 89.320 46.290 90.280 46.555 ;
        RECT 91.200 46.290 92.160 46.555 ;
        RECT 64.215 45.340 70.120 45.580 ;
        RECT 86.875 45.580 87.115 45.860 ;
        RECT 92.540 45.580 92.780 50.910 ;
        RECT 93.900 50.730 94.510 50.910 ;
        RECT 95.780 50.730 96.390 51.330 ;
        RECT 106.855 50.885 107.105 58.205 ;
        RECT 115.720 57.955 116.720 57.990 ;
        RECT 117.600 57.955 118.600 57.990 ;
        RECT 119.480 57.955 120.480 57.990 ;
        RECT 108.210 57.910 109.200 57.950 ;
        RECT 110.080 57.910 111.060 57.950 ;
        RECT 108.210 57.660 111.060 57.910 ;
        RECT 115.720 57.705 120.480 57.955 ;
        RECT 115.720 57.670 116.720 57.705 ;
        RECT 117.600 57.670 118.600 57.705 ;
        RECT 119.480 57.670 120.480 57.705 ;
        RECT 108.210 57.630 109.200 57.660 ;
        RECT 110.080 57.630 111.060 57.660 ;
        RECT 121.210 56.605 122.210 56.720 ;
        RECT 111.545 56.355 122.210 56.605 ;
        RECT 108.220 55.090 109.180 55.350 ;
        RECT 110.100 55.090 111.070 55.350 ;
        RECT 108.220 54.840 111.070 55.090 ;
        RECT 108.220 54.580 109.180 54.840 ;
        RECT 110.100 54.570 111.070 54.840 ;
        RECT 111.545 54.185 111.795 56.355 ;
        RECT 112.340 55.920 121.010 56.160 ;
        RECT 112.340 55.350 112.580 55.920 ;
        RECT 113.125 55.500 115.400 55.740 ;
        RECT 111.980 54.580 112.940 55.350 ;
        RECT 111.545 53.935 112.030 54.185 ;
        RECT 111.775 53.030 112.030 53.935 ;
        RECT 107.800 52.420 108.400 53.030 ;
        RECT 111.600 52.430 112.210 53.030 ;
        RECT 107.970 51.995 108.220 52.420 ;
        RECT 111.775 51.995 112.030 52.430 ;
        RECT 107.970 51.745 112.030 51.995 ;
        RECT 107.970 51.465 108.225 51.745 ;
        RECT 107.970 51.260 108.220 51.465 ;
        RECT 111.780 51.260 112.030 51.745 ;
        RECT 107.570 50.885 108.570 51.260 ;
        RECT 106.855 50.635 108.570 50.885 ;
        RECT 111.600 50.660 112.210 51.260 ;
        RECT 107.570 50.260 108.570 50.635 ;
        RECT 112.350 50.010 112.590 54.580 ;
        RECT 113.125 54.180 113.685 55.500 ;
        RECT 115.160 52.840 115.400 55.500 ;
        RECT 115.720 55.090 116.720 55.350 ;
        RECT 117.600 55.090 118.600 55.350 ;
        RECT 119.480 55.090 120.480 55.350 ;
        RECT 115.720 54.840 120.480 55.090 ;
        RECT 120.770 55.200 121.010 55.920 ;
        RECT 121.210 55.720 122.210 56.355 ;
        RECT 121.585 55.420 121.835 55.720 ;
        RECT 121.210 55.200 122.210 55.420 ;
        RECT 120.770 54.960 122.210 55.200 ;
        RECT 115.720 54.580 116.720 54.840 ;
        RECT 117.600 54.580 118.600 54.840 ;
        RECT 119.480 54.580 120.480 54.840 ;
        RECT 121.210 54.420 122.210 54.960 ;
        RECT 116.570 52.840 117.170 53.030 ;
        RECT 115.160 52.600 117.170 52.840 ;
        RECT 116.570 52.430 117.170 52.600 ;
        RECT 118.450 52.430 119.050 53.030 ;
        RECT 118.625 51.330 118.875 52.430 ;
        RECT 116.560 51.150 117.170 51.330 ;
        RECT 108.580 49.770 112.590 50.010 ;
        RECT 115.200 50.910 117.170 51.150 ;
        RECT 93.060 46.805 94.060 47.070 ;
        RECT 94.940 46.805 95.940 47.070 ;
        RECT 108.580 47.060 108.820 49.770 ;
        RECT 93.060 46.555 95.940 46.805 ;
        RECT 93.060 46.290 94.060 46.555 ;
        RECT 94.940 46.290 95.940 46.555 ;
        RECT 108.220 46.300 109.180 47.060 ;
        RECT 109.390 45.860 109.920 47.500 ;
        RECT 111.980 46.805 112.940 47.070 ;
        RECT 113.860 46.805 114.820 47.070 ;
        RECT 111.980 46.555 114.820 46.805 ;
        RECT 111.980 46.290 112.940 46.555 ;
        RECT 113.860 46.290 114.820 46.555 ;
        RECT 86.875 45.340 92.780 45.580 ;
        RECT 109.535 45.580 109.775 45.860 ;
        RECT 115.200 45.580 115.440 50.910 ;
        RECT 116.560 50.730 117.170 50.910 ;
        RECT 118.440 50.730 119.050 51.330 ;
        RECT 115.720 46.805 116.720 47.070 ;
        RECT 117.600 46.805 118.600 47.070 ;
        RECT 115.720 46.555 118.600 46.805 ;
        RECT 115.720 46.290 116.720 46.555 ;
        RECT 117.600 46.290 118.600 46.555 ;
        RECT 109.535 45.340 115.440 45.580 ;
        RECT 44.000 41.560 46.840 41.880 ;
        RECT 66.660 41.560 69.500 41.880 ;
        RECT 89.320 41.560 92.160 41.880 ;
        RECT 111.980 41.560 114.820 41.880 ;
      LAYER via2 ;
        RECT 51.530 176.590 51.810 176.870 ;
        RECT 57.510 165.030 57.790 165.310 ;
        RECT 59.350 173.870 59.630 174.150 ;
        RECT 67.170 165.030 67.450 165.310 ;
        RECT 70.850 177.270 71.130 177.550 ;
        RECT 73.150 171.830 73.430 172.110 ;
        RECT 73.150 163.670 73.430 163.950 ;
        RECT 82.810 174.550 83.090 174.830 ;
        RECT 82.810 169.110 83.090 169.390 ;
        RECT 89.250 177.270 89.530 177.550 ;
        RECT 86.030 174.550 86.310 174.830 ;
        RECT 82.350 165.710 82.630 165.990 ;
        RECT 87.410 171.150 87.690 171.430 ;
        RECT 86.950 169.110 87.230 169.390 ;
        RECT 91.090 171.150 91.370 171.430 ;
        RECT 91.550 169.110 91.830 169.390 ;
        RECT 95.230 173.190 95.510 173.470 ;
        RECT 96.610 177.270 96.890 177.550 ;
        RECT 99.370 165.710 99.650 165.990 ;
        RECT 108.570 176.590 108.850 176.870 ;
        RECT 104.890 171.830 105.170 172.110 ;
        RECT 109.490 172.510 109.770 172.790 ;
        RECT 105.810 163.670 106.090 163.950 ;
        RECT 104.890 160.270 105.170 160.550 ;
        RECT 109.490 171.150 109.770 171.430 ;
        RECT 112.250 169.110 112.530 169.390 ;
      LAYER met3 ;
        RECT 70.825 177.560 71.155 177.575 ;
        RECT 89.225 177.560 89.555 177.575 ;
        RECT 96.585 177.560 96.915 177.575 ;
        RECT 70.825 177.260 96.915 177.560 ;
        RECT 70.825 177.245 71.155 177.260 ;
        RECT 89.225 177.245 89.555 177.260 ;
        RECT 96.585 177.245 96.915 177.260 ;
        RECT 51.505 176.880 51.835 176.895 ;
        RECT 104.610 176.880 104.990 176.890 ;
        RECT 108.545 176.880 108.875 176.895 ;
        RECT 51.505 176.580 108.875 176.880 ;
        RECT 51.505 176.565 51.835 176.580 ;
        RECT 104.610 176.570 104.990 176.580 ;
        RECT 108.545 176.565 108.875 176.580 ;
        RECT 82.785 174.840 83.115 174.855 ;
        RECT 86.005 174.840 86.335 174.855 ;
        RECT 82.785 174.540 86.335 174.840 ;
        RECT 82.785 174.525 83.115 174.540 ;
        RECT 86.005 174.525 86.335 174.540 ;
        RECT 59.325 174.160 59.655 174.175 ;
        RECT 59.325 173.860 84.710 174.160 ;
        RECT 59.325 173.845 59.655 173.860 ;
        RECT 84.410 173.480 84.710 173.860 ;
        RECT 95.205 173.480 95.535 173.495 ;
        RECT 84.410 173.180 95.535 173.480 ;
        RECT 95.205 173.165 95.535 173.180 ;
        RECT 109.465 172.800 109.795 172.815 ;
        RECT 109.250 172.485 109.795 172.800 ;
        RECT 73.125 172.120 73.455 172.135 ;
        RECT 104.865 172.120 105.195 172.135 ;
        RECT 73.125 171.820 105.195 172.120 ;
        RECT 73.125 171.805 73.455 171.820 ;
        RECT 104.865 171.805 105.195 171.820 ;
        RECT 109.250 171.455 109.550 172.485 ;
        RECT 87.385 171.440 87.715 171.455 ;
        RECT 91.065 171.440 91.395 171.455 ;
        RECT 87.385 171.140 91.395 171.440 ;
        RECT 109.250 171.140 109.795 171.455 ;
        RECT 87.385 171.125 87.715 171.140 ;
        RECT 91.065 171.125 91.395 171.140 ;
        RECT 109.465 171.125 109.795 171.140 ;
        RECT 82.785 169.400 83.115 169.415 ;
        RECT 86.925 169.400 87.255 169.415 ;
        RECT 82.785 169.100 87.255 169.400 ;
        RECT 82.785 169.085 83.115 169.100 ;
        RECT 86.925 169.085 87.255 169.100 ;
        RECT 91.525 169.400 91.855 169.415 ;
        RECT 112.225 169.400 112.555 169.415 ;
        RECT 91.525 169.100 112.555 169.400 ;
        RECT 91.525 169.085 91.855 169.100 ;
        RECT 112.225 169.085 112.555 169.100 ;
        RECT 82.325 166.000 82.655 166.015 ;
        RECT 99.345 166.000 99.675 166.015 ;
        RECT 82.325 165.700 99.675 166.000 ;
        RECT 82.325 165.685 82.655 165.700 ;
        RECT 99.345 165.685 99.675 165.700 ;
        RECT 57.485 165.320 57.815 165.335 ;
        RECT 67.145 165.320 67.475 165.335 ;
        RECT 57.485 165.020 67.475 165.320 ;
        RECT 57.485 165.005 57.815 165.020 ;
        RECT 67.145 165.005 67.475 165.020 ;
        RECT 73.125 163.960 73.455 163.975 ;
        RECT 105.785 163.960 106.115 163.975 ;
        RECT 73.125 163.660 106.115 163.960 ;
        RECT 73.125 163.645 73.455 163.660 ;
        RECT 105.785 163.645 106.115 163.660 ;
        RECT 104.865 160.570 105.195 160.575 ;
        RECT 104.610 160.560 105.195 160.570 ;
        RECT 104.610 160.260 105.420 160.560 ;
        RECT 104.610 160.250 105.195 160.260 ;
        RECT 104.865 160.245 105.195 160.250 ;
      LAYER via3 ;
        RECT 104.640 176.570 104.960 176.890 ;
        RECT 104.640 160.250 104.960 160.570 ;
      LAYER met4 ;
        RECT 104.635 176.565 104.965 176.895 ;
        RECT 104.650 160.575 104.950 176.565 ;
        RECT 104.635 160.245 104.965 160.575 ;
  END
END tt_um_htfab_flash_adc
END LIBRARY

