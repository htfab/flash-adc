magic
tech sky130A
magscale 1 2
timestamp 1712769939
<< nwell >>
rect 850 -470 1610 -70
<< mvpdiff >>
rect 1090 -370 1116 -358
<< mvpsubdiff >>
rect 1494 -710 1536 -686
rect 1494 -776 1536 -752
<< mvnsubdiff >>
rect 1502 -194 1544 -170
rect 1502 -260 1544 -236
<< mvpsubdiffcont >>
rect 1494 -752 1536 -710
<< mvnsubdiffcont >>
rect 1502 -236 1544 -194
<< locali >>
rect 1502 -194 1544 -178
rect 1502 -252 1544 -236
rect 1494 -710 1536 -694
rect 1494 -768 1536 -752
<< viali >>
rect 1505 -231 1539 -197
rect 1498 -747 1532 -713
<< metal1 >>
rect 852 -55 1541 -17
rect 852 -70 890 -55
rect 690 -229 890 -70
rect 690 -267 968 -229
rect 690 -270 890 -267
rect 690 -475 890 -330
rect 1009 -450 1047 -89
rect 1167 -157 1205 -55
rect 1167 -195 1248 -157
rect 1087 -375 1163 -337
rect 978 -475 1047 -450
rect 690 -513 1047 -475
rect 690 -530 890 -513
rect 978 -544 1047 -513
rect 690 -654 890 -590
rect 690 -692 968 -654
rect 690 -759 890 -692
rect 690 -790 891 -759
rect 1009 -774 1047 -544
rect 1125 -473 1163 -375
rect 1289 -441 1327 -89
rect 1503 -185 1541 -55
rect 1499 -197 1545 -185
rect 1499 -231 1505 -197
rect 1539 -231 1545 -197
rect 1499 -243 1545 -231
rect 1368 -330 1406 -251
rect 1368 -375 1640 -330
rect 1257 -473 1327 -441
rect 1125 -511 1327 -473
rect 1125 -595 1163 -511
rect 1257 -556 1327 -511
rect 1087 -633 1163 -595
rect 1173 -702 1252 -664
rect 853 -811 891 -790
rect 1173 -811 1211 -702
rect 1289 -774 1327 -556
rect 1405 -530 1640 -375
rect 1405 -595 1443 -530
rect 1367 -633 1443 -595
rect 1492 -713 1538 -701
rect 1492 -747 1498 -713
rect 1532 -747 1538 -713
rect 1492 -759 1538 -747
rect 1496 -811 1533 -759
rect 853 -849 1533 -811
use cells/sky130_fd_pr__nfet_g5v0d10v5_VNEAGC  sky130_fd_pr__nfet_g5v0d10v5_VNEAGC_0 cells
timestamp 1712769939
transform 1 0 1028 0 1 -652
box -108 -138 108 138
use cells/sky130_fd_pr__nfet_g5v0d10v5_VNEAGC  sky130_fd_pr__nfet_g5v0d10v5_VNEAGC_2
timestamp 1712769939
transform 1 0 1308 0 1 -652
box -108 -138 108 138
use cells/sky130_fd_pr__pfet_g5v0d10v5_PC3LZ5  sky130_fd_pr__pfet_g5v0d10v5_PC3LZ5_0 cells
timestamp 1712769939
transform 1 0 1308 0 1 -270
box -174 -200 174 200
use cells/sky130_fd_pr__pfet_g5v0d10v5_PC3LZ5  sky130_fd_pr__pfet_g5v0d10v5_PC3LZ5_1
timestamp 1712769939
transform 1 0 1028 0 1 -270
box -174 -200 174 200
<< labels >>
flabel metal1 690 -790 890 -590 0 FreeSans 256 0 0 0 VSS
port 3 nsew
flabel metal1 690 -530 890 -330 0 FreeSans 256 0 0 0 IN
port 2 nsew
flabel metal1 1440 -530 1640 -330 0 FreeSans 256 0 0 0 OUT
port 1 nsew
flabel metal1 690 -270 890 -70 0 FreeSans 256 0 0 0 VDD
port 0 nsew
<< end >>
