magic
tech sky130A
magscale 1 2
timestamp 1713023969
<< metal1 >>
rect 1258 1278 1328 1284
rect 1258 840 1328 846
rect 1258 378 1328 384
rect 1258 -60 1328 -54
rect 1258 -280 1328 -274
rect 5404 -320 5604 -312
rect 5404 -504 5412 -320
rect 5596 -504 5604 -320
rect 5404 -512 5604 -504
rect 1258 -718 1328 -712
rect 4906 -969 4972 -888
rect 5026 -969 5092 -888
rect 5146 -969 5212 -888
rect 5266 -969 5332 -888
rect 5547 -969 5597 -512
rect 4906 -1019 5597 -969
rect 4906 -1100 4972 -1019
rect 5026 -1100 5092 -1019
rect 5146 -1100 5212 -1019
rect 5266 -1100 5332 -1019
rect 1726 -1158 1864 -1144
rect 1258 -1180 1328 -1174
rect 1506 -1270 1512 -1218
rect 1564 -1225 1570 -1218
rect 1726 -1225 1742 -1158
rect 1564 -1263 1742 -1225
rect 1564 -1270 1570 -1263
rect 1726 -1330 1742 -1263
rect 1850 -1330 1864 -1158
rect 1726 -1344 1864 -1330
rect 1258 -1618 1328 -1612
<< via1 >>
rect 1258 846 1328 1278
rect 1258 -54 1328 378
rect 1258 -712 1328 -280
rect 5412 -504 5596 -320
rect 1258 -1612 1328 -1180
rect 1512 -1270 1564 -1218
rect 1742 -1330 1850 -1158
<< metal2 >>
rect 1268 1284 1318 1538
rect 1258 1278 1328 1284
rect 1258 840 1328 846
rect 1258 378 1328 384
rect 1258 -60 1328 -54
rect 1268 -141 1318 -60
rect 1268 -191 1563 -141
rect 1268 -274 1318 -191
rect 1258 -280 1328 -274
rect 1258 -718 1328 -712
rect 1258 -1180 1328 -1174
rect 1513 -1212 1563 -191
rect 1608 -963 1658 1538
rect 5404 -320 5604 -312
rect 5404 -504 5412 -320
rect 5596 -504 5604 -320
rect 5404 -512 5604 -504
rect 1726 -640 1926 -630
rect 1726 -820 1736 -640
rect 1916 -820 1926 -640
rect 1726 -830 1926 -820
rect 1608 -1013 1851 -963
rect 1512 -1218 1564 -1212
rect 1512 -1276 1564 -1270
rect 1258 -1618 1328 -1612
rect 1268 -1858 1318 -1618
rect 1608 -1858 1658 -1013
rect 1726 -1668 1926 -1658
rect 1726 -1848 1736 -1668
rect 1916 -1848 1926 -1668
rect 1726 -1858 1926 -1848
<< via2 >>
rect 1736 -820 1916 -640
rect 1736 -1848 1916 -1668
<< metal3 >>
rect 1092 306 5604 506
rect 1726 -640 1926 306
rect 1726 -820 1736 -640
rect 1916 -820 1926 -640
rect 1726 -830 1926 -820
rect 1092 -1344 5604 -1144
rect 1726 -1668 1926 -1344
rect 1726 -1848 1736 -1668
rect 1916 -1848 1926 -1668
rect 1726 -1858 1926 -1848
use comparator  comparator_0
timestamp 1713023969
transform 1 0 1356 0 1 -264
box 370 -1594 4248 1802
use cells/sky130_fd_pr__res_xhigh_po_0p35_29QZGQ  sky130_fd_pr__res_xhigh_po_0p35_29QZGQ_0 cells
timestamp 1713023969
transform 1 0 1293 0 1 612
box -201 -832 201 832
use cells/sky130_fd_pr__res_xhigh_po_0p35_29QZGQ  sky130_fd_pr__res_xhigh_po_0p35_29QZGQ_1
timestamp 1713023969
transform 1 0 1293 0 1 -946
box -201 -832 201 832
<< labels >>
flabel metal2 1608 -1858 1658 -1658 0 FreeSans 256 0 0 0 IN
port 2 nsew
flabel metal2 1608 1338 1658 1538 0 FreeSans 256 0 0 0 IN
port 2 nsew
flabel metal2 5404 -512 5604 -312 0 FreeSans 256 0 0 0 OUT
port 3 nsew
flabel metal3 1092 306 5604 506 0 FreeSans 256 0 0 0 VDD
port 1 nsew
flabel metal3 1092 -1344 5604 -1144 0 FreeSans 256 0 0 0 VSS
port 4 nsew
flabel metal1 4912 -1094 4966 -894 0 FreeSans 256 0 0 0 OUT
port 1 nsew
flabel metal1 5032 -1094 5086 -894 0 FreeSans 256 0 0 0 OUT
port 1 nsew
flabel metal1 5152 -1094 5206 -894 0 FreeSans 256 0 0 0 OUT
port 1 nsew
flabel metal1 5272 -1094 5326 -894 0 FreeSans 256 0 0 0 OUT
port 1 nsew
flabel metal2 1268 -1858 1318 -1658 0 FreeSans 256 0 0 0 REF1
port 5 nsew
flabel metal2 1268 1338 1318 1538 0 FreeSans 256 0 0 0 REF2
port 0 nsew
<< end >>
